
--------------------------------------------------------------------------------
-- End of file
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--       ------------      Project : bit_ser_adder
--    ,' GoodLuck ,'      RCSfile: ha.vhd,v  
--   '-----------'     Author: DR \*
--
--  Revision: 1.1  
--  Date: 1999.12.31
--  State: Exp  
--  Locker:   
--------------------------------------------------------------------------------
--
-- Description : Half adder
--
--
--------------------------------------------------------------------------------
--
--  Source: ./git/COMMON/IPs/NLWARE/DSP/bit_ser_adder/vhdl/rtl/ha.vhd,v  
--  Log: ha.vhd,v  
-- Revision 1.1  2003/04/18 07:07:56  rrich
-- Initial revision
--
--
--
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Library
--------------------------------------------------------------------------------
library IEEE; 
use IEEE.STD_LOGIC_1164.ALL;

--------------------------------------------------------------------------------
-- Entity
--------------------------------------------------------------------------------
entity ha is
  
  port (
    x : in  std_logic;
    y : in  std_logic;
    c : out std_logic;
    s : out std_logic);
    
end ha;
