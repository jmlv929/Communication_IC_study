
/*Vx2, V2.1.5
Released 2006-10-10
Checked out from CVS as $Header: //acds/rel/13.0sp1/ip/infrastructure/tools/lib/ToolVersion.pm#1 $
*/// vx_version verilog
// vx_version
/*
***********************************************************
title:   encoding_lut.vx
desc:    Encoder Look Up Table
author:  Enang Akan, eakan@altera.com
         www.altera.com   (c) 2002 Altera OTC Inc.
         tel: (613) 591-6700  fax: (613) 591-6831
***********************************************************
*/
module  b8tob10_encoding_lut (
reset_n,
clk,
rdaddress_a,
q_a);

// Ports and local variables. 
// '_F' indicates an auxiliary variable for flip-flops
// '_S' indicates an auxiliary variable for combinational signals
// '_W' indicates a VX2-created wire
input reset_n;
input clk;
input[7:0] rdaddress_a;
output[15:0] q_a;
wire  reset_n ;
wire  clk ;
wire  [7:0] rdaddress_a  ;
reg  [15:0] q_a, _Fq_a  ;
reg  [15:0] q_pre1_a, _Sq_pre1_a  ;

always @( * )  begin
// initialize flip-flop and combinational regs
    _Fq_a = q_a;
    _Sq_pre1_a = 0;

// mainline code
    begin // *** put code block here *** 

        case (rdaddress_a)
            0:
                _Sq_pre1_a = 16'b0001110010111001;
            1:
                _Sq_pre1_a = 16'b0001110010101110;
            2:
                _Sq_pre1_a = 16'b0001110010101101;
            3:
                _Sq_pre1_a = 16'b0001001101100011;
            4:
                _Sq_pre1_a = 16'b0001110010101011;
            5:
                _Sq_pre1_a = 16'b0001001101100101;
            6:
                _Sq_pre1_a = 16'b0001001101100110;
            7:
                _Sq_pre1_a = 16'b0001101101000111;
            8:
                _Sq_pre1_a = 16'b0001110010100111;
            9:
                _Sq_pre1_a = 16'b0001001101101001;
            10:
                _Sq_pre1_a = 16'b0001001101101010;
            11:
                _Sq_pre1_a = 16'b0001001101001011;
            12:
                _Sq_pre1_a = 16'b0001001101101100;
            13:
                _Sq_pre1_a = 16'b0001001101001101;
            14:
                _Sq_pre1_a = 16'b0001001101001110;
            15:
                _Sq_pre1_a = 16'b0001110010111010;
            16:
                _Sq_pre1_a = 16'b0001110010110110;
            17:
                _Sq_pre1_a = 16'b0001001101110001;
            18:
                _Sq_pre1_a = 16'b0001001101110010;
            19:
                _Sq_pre1_a = 16'b0001001101010011;
            20:
                _Sq_pre1_a = 16'b0001001101110100;
            21:
                _Sq_pre1_a = 16'b0001001101010101;
            22:
                _Sq_pre1_a = 16'b0001001101010110;
            23:
                _Sq_pre1_a = 16'b0001110010010111;
            24:
                _Sq_pre1_a = 16'b0001110010110011;
            25:
                _Sq_pre1_a = 16'b0001001101011001;
            26:
                _Sq_pre1_a = 16'b0001001101011010;
            27:
                _Sq_pre1_a = 16'b0001110010011011;
            28:
                _Sq_pre1_a = 16'b1101001101011100;
            29:
                _Sq_pre1_a = 16'b0001110010011101;
            30:
                _Sq_pre1_a = 16'b0001110010011110;
            31:
                _Sq_pre1_a = 16'b0001110010110101;
            32:
                _Sq_pre1_a = 16'b0000101001111001;
            33:
                _Sq_pre1_a = 16'b0000101001101110;
            34:
                _Sq_pre1_a = 16'b0000101001101101;
            35:
                _Sq_pre1_a = 16'b0000011001100011;
            36:
                _Sq_pre1_a = 16'b0000101001101011;
            37:
                _Sq_pre1_a = 16'b0000011001100101;
            38:
                _Sq_pre1_a = 16'b0000011001100110;
            39:
                _Sq_pre1_a = 16'b0000111001000111;
            40:
                _Sq_pre1_a = 16'b0000101001100111;
            41:
                _Sq_pre1_a = 16'b0000011001101001;
            42:
                _Sq_pre1_a = 16'b0000011001101010;
            43:
                _Sq_pre1_a = 16'b0000011001001011;
            44:
                _Sq_pre1_a = 16'b0000011001101100;
            45:
                _Sq_pre1_a = 16'b0000011001001101;
            46:
                _Sq_pre1_a = 16'b0000011001001110;
            47:
                _Sq_pre1_a = 16'b0000101001111010;
            48:
                _Sq_pre1_a = 16'b0000101001110110;
            49:
                _Sq_pre1_a = 16'b0000011001110001;
            50:
                _Sq_pre1_a = 16'b0000011001110010;
            51:
                _Sq_pre1_a = 16'b0000011001010011;
            52:
                _Sq_pre1_a = 16'b0000011001110100;
            53:
                _Sq_pre1_a = 16'b0000011001010101;
            54:
                _Sq_pre1_a = 16'b0000011001010110;
            55:
                _Sq_pre1_a = 16'b0000101001010111;
            56:
                _Sq_pre1_a = 16'b0000101001110011;
            57:
                _Sq_pre1_a = 16'b0000011001011001;
            58:
                _Sq_pre1_a = 16'b0000011001011010;
            59:
                _Sq_pre1_a = 16'b0000101001011011;
            60:
                _Sq_pre1_a = 16'b1000011001011100;
            61:
                _Sq_pre1_a = 16'b0000101001011101;
            62:
                _Sq_pre1_a = 16'b0000101001011110;
            63:
                _Sq_pre1_a = 16'b0000101001110101;
            64:
                _Sq_pre1_a = 16'b0000101010111001;
            65:
                _Sq_pre1_a = 16'b0000101010101110;
            66:
                _Sq_pre1_a = 16'b0000101010101101;
            67:
                _Sq_pre1_a = 16'b0000011010100011;
            68:
                _Sq_pre1_a = 16'b0000101010101011;
            69:
                _Sq_pre1_a = 16'b0000011010100101;
            70:
                _Sq_pre1_a = 16'b0000011010100110;
            71:
                _Sq_pre1_a = 16'b0000111010000111;
            72:
                _Sq_pre1_a = 16'b0000101010100111;
            73:
                _Sq_pre1_a = 16'b0000011010101001;
            74:
                _Sq_pre1_a = 16'b0000011010101010;
            75:
                _Sq_pre1_a = 16'b0000011010001011;
            76:
                _Sq_pre1_a = 16'b0000011010101100;
            77:
                _Sq_pre1_a = 16'b0000011010001101;
            78:
                _Sq_pre1_a = 16'b0000011010001110;
            79:
                _Sq_pre1_a = 16'b0000101010111010;
            80:
                _Sq_pre1_a = 16'b0000101010110110;
            81:
                _Sq_pre1_a = 16'b0000011010110001;
            82:
                _Sq_pre1_a = 16'b0000011010110010;
            83:
                _Sq_pre1_a = 16'b0000011010010011;
            84:
                _Sq_pre1_a = 16'b0000011010110100;
            85:
                _Sq_pre1_a = 16'b0000011010010101;
            86:
                _Sq_pre1_a = 16'b0000011010010110;
            87:
                _Sq_pre1_a = 16'b0000101010010111;
            88:
                _Sq_pre1_a = 16'b0000101010110011;
            89:
                _Sq_pre1_a = 16'b0000011010011001;
            90:
                _Sq_pre1_a = 16'b0000011010011010;
            91:
                _Sq_pre1_a = 16'b0000101010011011;
            92:
                _Sq_pre1_a = 16'b1000011010011100;
            93:
                _Sq_pre1_a = 16'b0000101010011101;
            94:
                _Sq_pre1_a = 16'b0000101010011110;
            95:
                _Sq_pre1_a = 16'b0000101010110101;
            96:
                _Sq_pre1_a = 16'b0001101100111001;
            97:
                _Sq_pre1_a = 16'b0001101100101110;
            98:
                _Sq_pre1_a = 16'b0001101100101101;
            99:
                _Sq_pre1_a = 16'b0001010011100011;
            100:
                _Sq_pre1_a = 16'b0001101100101011;
            101:
                _Sq_pre1_a = 16'b0001010011100101;
            102:
                _Sq_pre1_a = 16'b0001010011100110;
            103:
                _Sq_pre1_a = 16'b0001110011000111;
            104:
                _Sq_pre1_a = 16'b0001101100100111;
            105:
                _Sq_pre1_a = 16'b0001010011101001;
            106:
                _Sq_pre1_a = 16'b0001010011101010;
            107:
                _Sq_pre1_a = 16'b0001010011001011;
            108:
                _Sq_pre1_a = 16'b0001010011101100;
            109:
                _Sq_pre1_a = 16'b0001010011001101;
            110:
                _Sq_pre1_a = 16'b0001010011001110;
            111:
                _Sq_pre1_a = 16'b0001101100111010;
            112:
                _Sq_pre1_a = 16'b0001101100110110;
            113:
                _Sq_pre1_a = 16'b0001010011110001;
            114:
                _Sq_pre1_a = 16'b0001010011110010;
            115:
                _Sq_pre1_a = 16'b0001010011010011;
            116:
                _Sq_pre1_a = 16'b0001010011110100;
            117:
                _Sq_pre1_a = 16'b0001010011010101;
            118:
                _Sq_pre1_a = 16'b0001010011010110;
            119:
                _Sq_pre1_a = 16'b0001101100010111;
            120:
                _Sq_pre1_a = 16'b0001101100110011;
            121:
                _Sq_pre1_a = 16'b0001010011011001;
            122:
                _Sq_pre1_a = 16'b0001010011011010;
            123:
                _Sq_pre1_a = 16'b0001101100011011;
            124:
                _Sq_pre1_a = 16'b1001010011011100;
            125:
                _Sq_pre1_a = 16'b0001101100011101;
            126:
                _Sq_pre1_a = 16'b0001101100011110;
            127:
                _Sq_pre1_a = 16'b0001101100110101;
            128:
                _Sq_pre1_a = 16'b0001110100111001;
            129:
                _Sq_pre1_a = 16'b0001110100101110;
            130:
                _Sq_pre1_a = 16'b0001110100101101;
            131:
                _Sq_pre1_a = 16'b0001001011100011;
            132:
                _Sq_pre1_a = 16'b0001110100101011;
            133:
                _Sq_pre1_a = 16'b0001001011100101;
            134:
                _Sq_pre1_a = 16'b0001001011100110;
            135:
                _Sq_pre1_a = 16'b0001101011000111;
            136:
                _Sq_pre1_a = 16'b0001110100100111;
            137:
                _Sq_pre1_a = 16'b0001001011101001;
            138:
                _Sq_pre1_a = 16'b0001001011101010;
            139:
                _Sq_pre1_a = 16'b0001001011001011;
            140:
                _Sq_pre1_a = 16'b0001001011101100;
            141:
                _Sq_pre1_a = 16'b0001001011001101;
            142:
                _Sq_pre1_a = 16'b0001001011001110;
            143:
                _Sq_pre1_a = 16'b0001110100111010;
            144:
                _Sq_pre1_a = 16'b0001110100110110;
            145:
                _Sq_pre1_a = 16'b0001001011110001;
            146:
                _Sq_pre1_a = 16'b0001001011110010;
            147:
                _Sq_pre1_a = 16'b0001001011010011;
            148:
                _Sq_pre1_a = 16'b0001001011110100;
            149:
                _Sq_pre1_a = 16'b0001001011010101;
            150:
                _Sq_pre1_a = 16'b0001001011010110;
            151:
                _Sq_pre1_a = 16'b0001110100010111;
            152:
                _Sq_pre1_a = 16'b0001110100110011;
            153:
                _Sq_pre1_a = 16'b0001001011011001;
            154:
                _Sq_pre1_a = 16'b0001001011011010;
            155:
                _Sq_pre1_a = 16'b0001110100011011;
            156:
                _Sq_pre1_a = 16'b1101001011011100;
            157:
                _Sq_pre1_a = 16'b0001110100011101;
            158:
                _Sq_pre1_a = 16'b0001110100011110;
            159:
                _Sq_pre1_a = 16'b0001110100110101;
            160:
                _Sq_pre1_a = 16'b0000100101111001;
            161:
                _Sq_pre1_a = 16'b0000100101101110;
            162:
                _Sq_pre1_a = 16'b0000100101101101;
            163:
                _Sq_pre1_a = 16'b0000010101100011;
            164:
                _Sq_pre1_a = 16'b0000100101101011;
            165:
                _Sq_pre1_a = 16'b0000010101100101;
            166:
                _Sq_pre1_a = 16'b0000010101100110;
            167:
                _Sq_pre1_a = 16'b0000110101000111;
            168:
                _Sq_pre1_a = 16'b0000100101100111;
            169:
                _Sq_pre1_a = 16'b0000010101101001;
            170:
                _Sq_pre1_a = 16'b0000010101101010;
            171:
                _Sq_pre1_a = 16'b0000010101001011;
            172:
                _Sq_pre1_a = 16'b0000010101101100;
            173:
                _Sq_pre1_a = 16'b0000010101001101;
            174:
                _Sq_pre1_a = 16'b0000010101001110;
            175:
                _Sq_pre1_a = 16'b0000100101111010;
            176:
                _Sq_pre1_a = 16'b0000100101110110;
            177:
                _Sq_pre1_a = 16'b0000010101110001;
            178:
                _Sq_pre1_a = 16'b0000010101110010;
            179:
                _Sq_pre1_a = 16'b0000010101010011;
            180:
                _Sq_pre1_a = 16'b0000010101110100;
            181:
                _Sq_pre1_a = 16'b0000010101010101;
            182:
                _Sq_pre1_a = 16'b0000010101010110;
            183:
                _Sq_pre1_a = 16'b0000100101010111;
            184:
                _Sq_pre1_a = 16'b0000100101110011;
            185:
                _Sq_pre1_a = 16'b0000010101011001;
            186:
                _Sq_pre1_a = 16'b0000010101011010;
            187:
                _Sq_pre1_a = 16'b0000100101011011;
            188:
                _Sq_pre1_a = 16'b1000010101011100;
            189:
                _Sq_pre1_a = 16'b0000100101011101;
            190:
                _Sq_pre1_a = 16'b0000100101011110;
            191:
                _Sq_pre1_a = 16'b0000100101110101;
            192:
                _Sq_pre1_a = 16'b0000100110111001;
            193:
                _Sq_pre1_a = 16'b0000100110101110;
            194:
                _Sq_pre1_a = 16'b0000100110101101;
            195:
                _Sq_pre1_a = 16'b0000010110100011;
            196:
                _Sq_pre1_a = 16'b0000100110101011;
            197:
                _Sq_pre1_a = 16'b0000010110100101;
            198:
                _Sq_pre1_a = 16'b0000010110100110;
            199:
                _Sq_pre1_a = 16'b0000110110000111;
            200:
                _Sq_pre1_a = 16'b0000100110100111;
            201:
                _Sq_pre1_a = 16'b0000010110101001;
            202:
                _Sq_pre1_a = 16'b0000010110101010;
            203:
                _Sq_pre1_a = 16'b0000010110001011;
            204:
                _Sq_pre1_a = 16'b0000010110101100;
            205:
                _Sq_pre1_a = 16'b0000010110001101;
            206:
                _Sq_pre1_a = 16'b0000010110001110;
            207:
                _Sq_pre1_a = 16'b0000100110111010;
            208:
                _Sq_pre1_a = 16'b0000100110110110;
            209:
                _Sq_pre1_a = 16'b0000010110110001;
            210:
                _Sq_pre1_a = 16'b0000010110110010;
            211:
                _Sq_pre1_a = 16'b0000010110010011;
            212:
                _Sq_pre1_a = 16'b0000010110110100;
            213:
                _Sq_pre1_a = 16'b0000010110010101;
            214:
                _Sq_pre1_a = 16'b0000010110010110;
            215:
                _Sq_pre1_a = 16'b0000100110010111;
            216:
                _Sq_pre1_a = 16'b0000100110110011;
            217:
                _Sq_pre1_a = 16'b0000010110011001;
            218:
                _Sq_pre1_a = 16'b0000010110011010;
            219:
                _Sq_pre1_a = 16'b0000100110011011;
            220:
                _Sq_pre1_a = 16'b1000010110011100;
            221:
                _Sq_pre1_a = 16'b0000100110011101;
            222:
                _Sq_pre1_a = 16'b0000100110011110;
            223:
                _Sq_pre1_a = 16'b0000100110110101;
            224:
                _Sq_pre1_a = 16'b0001111000111001;
            225:
                _Sq_pre1_a = 16'b0001111000101110;
            226:
                _Sq_pre1_a = 16'b0001111000101101;
            227:
                _Sq_pre1_a = 16'b0001000111100011;
            228:
                _Sq_pre1_a = 16'b0001111000101011;
            229:
                _Sq_pre1_a = 16'b0001000111100101;
            230:
                _Sq_pre1_a = 16'b0001000111100110;
            231:
                _Sq_pre1_a = 16'b0001100111000111;
            232:
                _Sq_pre1_a = 16'b0001111000100111;
            233:
                _Sq_pre1_a = 16'b0001000111101001;
            234:
                _Sq_pre1_a = 16'b0001000111101010;
            235:
                _Sq_pre1_a = 16'b0010000111001011;
            236:
                _Sq_pre1_a = 16'b0001000111101100;
            237:
                _Sq_pre1_a = 16'b0010000111001101;
            238:
                _Sq_pre1_a = 16'b0010000111001110;
            239:
                _Sq_pre1_a = 16'b0001111000111010;
            240:
                _Sq_pre1_a = 16'b0001111000110110;
            241:
                _Sq_pre1_a = 16'b0010001110110001;
            242:
                _Sq_pre1_a = 16'b0010001110110010;
            243:
                _Sq_pre1_a = 16'b0001000111010011;
            244:
                _Sq_pre1_a = 16'b0010001110110100;
            245:
                _Sq_pre1_a = 16'b0001000111010101;
            246:
                _Sq_pre1_a = 16'b0001000111010110;
            247:
                _Sq_pre1_a = 16'b1101111000010111;
            248:
                _Sq_pre1_a = 16'b0001111000110011;
            249:
                _Sq_pre1_a = 16'b0001000111011001;
            250:
                _Sq_pre1_a = 16'b0001000111011010;
            251:
                _Sq_pre1_a = 16'b1101111000011011;
            252:
                _Sq_pre1_a = 16'b1101000111011100;
            253:
                _Sq_pre1_a = 16'b1101111000011101;
            254:
                _Sq_pre1_a = 16'b1101111000011110;
            255:
                _Sq_pre1_a = 16'b1101111000110101;
        endcase
        _Fq_a = q_pre1_a;
    end 


// update regs for combinational signals
// The non-blocking assignment causes the always block to 
// re-stimulate if the signal has changed
    q_pre1_a <= _Sq_pre1_a;
end
always @(posedge clk or negedge reset_n) begin
    if (!reset_n) begin
        q_a<=0;
    end else begin
        q_a<=_Fq_a;
    end
end
endmodule
