

--------------------------------------------------------------------------------
-- Architecture
--------------------------------------------------------------------------------
architecture RTL of key_mixing_sbox is

  ------------------------------------------------------------------------------
  -- Types
  ------------------------------------------------------------------------------
  type SBOX_ARRAY_TYPE is array(0 to 255) of std_logic_vector(15 downto 0);

  ------------------------------------------------------------------------------
  -- Constants
  ------------------------------------------------------------------------------
  constant SBOX_TABLE_CT : SBOX_ARRAY_TYPE := (
    "1100011010100101", "1111100010000100", "1110111010011001", "1111011010001101", "1111111100001101", "1101011010111101", "1101111010110001", "1001000101010100",
    "0110000001010000", "0000001000000011", "1100111010101001", "0101011001111101", "1110011100011001", "1011010101100010", "0100110111100110", "1110110010011010",
    "1000111101000101", "0001111110011101", "1000100101000000", "1111101010000111", "1110111100010101", "1011001011101011", "1000111011001001", "1111101100001011",
    "0100000111101100", "1011001101100111", "0101111111111101", "0100010111101010", "0010001110111111", "0101001111110111", "1110010010010110", "1001101101011011",
    "0111010111000010", "1110000100011100", "0011110110101110", "0100110001101010", "0110110001011010", "0111111001000001", "1111010100000010", "1000001101001111",
    "0110100001011100", "0101000111110100", "1101000100110100", "1111100100001000", "1110001010010011", "1010101101110011", "0110001001010011", "0010101000111111",
    "0000100000001100", "1001010101010010", "0100011001100101", "1001110101011110", "0011000000101000", "0011011110100001", "0000101000001111", "0010111110110101",
    "0000111000001001", "0010010000110110", "0001101110011011", "1101111100111101", "1100110100100110", "0100111001101001", "0111111111001101", "1110101010011111",
    "0001001000011011", "0001110110011110", "0101100001110100", "0011010000101110", "0011011000101101", "1101110010110010", "1011010011101110", "0101101111111011",
    "1010010011110110", "0111011001001101", "1011011101100001", "0111110111001110", "0101001001111011", "1101110100111110", "0101111001110001", "0001001110010111",
    "1010011011110101", "1011100101101000", "0000000000000000", "1100000100101100", "0100000001100000", "1110001100011111", "0111100111001000", "1011011011101101",
    "1101010010111110", "1000110101000110", "0110011111011001", "0111001001001011", "1001010011011110", "1001100011010100", "1011000011101000", "1000010101001010",
    "1011101101101011", "1100010100101010", "0100111111100101", "1110110100010110", "1000011011000101", "1001101011010111", "0110011001010101", "0001000110010100",
    "1000101011001111", "1110100100010000", "0000010000000110", "1111111010000001", "1010000011110000", "0111100001000100", "0010010110111010", "0100101111100011",
    "1010001011110011", "0101110111111110", "1000000011000000", "0000010110001010", "0011111110101101", "0010000110111100", "0111000001001000", "1111000100000100",
    "0110001111011111", "0111011111000001", "1010111101110101", "0100001001100011", "0010000000110000", "1110010100011010", "1111110100001110", "1011111101101101",
    "1000000101001100", "0001100000010100", "0010011000110101", "1100001100101111", "1011111011100001", "0011010110100010", "1000100011001100", "0010111000111001",
    "1001001101010111", "0101010111110010", "1111110010000010", "0111101001000111", "1100100010101100", "1011101011100111", "0011001000101011", "1110011010010101",
    "1100000010100000", "0001100110011000", "1001111011010001", "1010001101111111", "0100010001100110", "0101010001111110", "0011101110101011", "0000101110000011",
    "1000110011001010", "1100011100101001", "0110101111010011", "0010100000111100", "1010011101111001", "1011110011100010", "0001011000011101", "1010110101110110",
    "1101101100111011", "0110010001010110", "0111010001001110", "0001010000011110", "1001001011011011", "0000110000001010", "0100100001101100", "1011100011100100",
    "1001111101011101", "1011110101101110", "0100001111101111", "1100010010100110", "0011100110101000", "0011000110100100", "1101001100110111", "1111001010001011",
    "1101010100110010", "1000101101000011", "0110111001011001", "1101101010110111", "0000000110001100", "1011000101100100", "1001110011010010", "0100100111100000",
    "1101100010110100", "1010110011111010", "1111001100000111", "1100111100100101", "1100101010101111", "1111010010001110", "0100011111101001", "0001000000011000",
    "0110111111010101", "1111000010001000", "0100101001101111", "0101110001110010", "0011100000100100", "0101011111110001", "0111001111000111", "1001011101010001",
    "1100101100100011", "1010000101111100", "1110100010011100", "0011111000100001", "1001011011011101", "0110000111011100", "0000110110000110", "0000111110000101",
    "1110000010010000", "0111110001000010", "0111000111000100", "1100110010101010", "1001000011011000", "0000011000000101", "1111011100000001", "0001110000010010",
    "1100001010100011", "0110101001011111", "1010111011111001", "0110100111010000", "0001011110010001", "1001100101011000", "0011101000100111", "0010011110111001",
    "1101100100111000", "1110101100010011", "0010101110110011", "0010001000110011", "1101001010111011", "1010100101110000", "0000011110001001", "0011001110100111",
    "0010110110110110", "0011110000100010", "0001010110010010", "1100100100100000", "1000011101001001", "1010101011111111", "0101000001111000", "1010010101111010",
    "0000001110001111", "0101100111111000", "0000100110000000", "0001101000010111", "0110010111011010", "1101011100110001", "1000010011000110", "1101000010111000",
    "1000001011000011", "0010100110110000", "0101101001110111", "0001111000010001", "0111101111001011", "1010100011111100", "0110110111010110", "0010110000111010");

  ------------------------------------------------------------------------------
  -- Signals
  ------------------------------------------------------------------------------
  signal sbox_data0 : std_logic_vector(15 downto 0);
  signal sbox_data1 : std_logic_vector(15 downto 0);
  
--------------------------------------------------------------------------------
-- Architecture Body
--------------------------------------------------------------------------------
begin
  sbox_data0 <= SBOX_TABLE_CT(conv_integer(sbox_addr(7 downto 0)));
  
  sbox1_pr: process(sbox_addr)
    variable sbox1_v : std_logic_vector(15 downto 0);
  begin
    sbox1_v := SBOX_TABLE_CT(conv_integer(sbox_addr(15 downto 8)));
    sbox_data1 <= sbox1_v(7 downto 0) & sbox1_v(15 downto 8);
  end process sbox1_pr;
  
  sbox_data <= sbox_data0 xor sbox_data1;

end RTL;
