// -------------------------------------------------------------
// HDL Code Generation Options:
//
// ResetType: Synchronous
// FIRAdderStyle: tree
// ResetInputPort: syn_rst
// TargetDirectory: E:\�ٶ���ͬ����\�鼮\���\������
// Name: fir_da
// RemoveResetFrom: ShiftRegister
// DALUTPartition: 5
// DARadix: 256
// TargetLanguage: Verilog
// TestBenchStimulus: impulse step ramp chirp noise 
//
// Filter Settings:
//
// Discrete-Time FIR Filter (real)
// -------------------------------
// Filter Structure  : Direct-Form FIR
// Filter Length     : 5
// Stable            : Yes
// Linear Phase      : Yes (Type 1)
// Arithmetic        : fixed
// Numerator         : s16,19 -> [-6.250000e-02 6.250000e-02)
// Input             : s8,7 -> [-1 1)
// Filter Internals  : Specify Precision
//   Output          : s8,7 -> [-1 1)
//   Product         : s31,31 -> [-5.000000e-01 5.000000e-01)
//   Accumulator     : s33,31 -> [-2 2)
//   Round Mode      : convergent
//   Overflow Mode   : wrap
// -------------------------------------------------------------
`timescale 1 ns / 1 ns 

module filter_tb;

// Function definitions
   function signed [7:0] abs;
   input signed [7:0] arg;
   begin
     abs = arg > 0 ? arg : -arg;
   end
   endfunction // function abs

  task filter_in_data_log_task; 
    input          clk;
    input          reset;
    input          rdenb;
    inout  [11:0]  addr;
    output         done;
  begin

    // Counter to generate the address
    if (reset == 1) 
      addr = 0;
    else begin
      if (rdenb == 1) begin
        if (addr == 3106)
          addr = addr; 
        else
          addr =  addr + 1; 
      end
    end

    // Done Signal generation.
    if (reset == 1)
      done = 0; 
    else if (addr == 3106)
      done = 1; 
    else
      done = 0; 

  end
  endtask // filter_in_data_log_task

  task filter_out_task; 
    input          clk;
    input          reset;
    input          rdenb;
    inout  [11:0]  addr;
    output         done;
  begin

    // Counter to generate the address
    if (reset == 1) 
      addr = 0;
    else begin
      if (rdenb == 1) begin
        if (addr == 3106)
          addr = addr; 
        else
          addr = #1  addr + 1; 
      end
    end

    // Done Signal generation.
    if (reset == 1)
      done = 0; 
    else if (addr == 3106)
      done = 1; 
    else
      done = 0; 

  end
  endtask // filter_out_task

 // Constants
 parameter clk_high                         = 5;
 parameter clk_low                          = 5;
 parameter clk_period                       = 10;
 parameter clk_hold                         = 2;
// -------------------------------------------------------------
//
// Module: filter_tb_data
// Generated by MATLAB(R) 8.3 and the Filter Design HDL Coder 2.9.5.
// Generated on: 2015-01-02 09:32:22
// -------------------------------------------------------------

  reg  signed [7:0] filter_in_data_log_force [0:3106];
  reg  signed [7:0] filter_out_expected [0:3106];


// **************************************
  initial //Input & Output data
  begin

  // Input data for filter_in_data_log
  filter_in_data_log_force[   0] <= 8'h7f;
  filter_in_data_log_force[   1] <= 8'h00;
  filter_in_data_log_force[   2] <= 8'h00;
  filter_in_data_log_force[   3] <= 8'h00;
  filter_in_data_log_force[   4] <= 8'h00;
  filter_in_data_log_force[   5] <= 8'h00;
  filter_in_data_log_force[   6] <= 8'h00;
  filter_in_data_log_force[   7] <= 8'h00;
  filter_in_data_log_force[   8] <= 8'h00;
  filter_in_data_log_force[   9] <= 8'h00;
  filter_in_data_log_force[  10] <= 8'h00;
  filter_in_data_log_force[  11] <= 8'h7f;
  filter_in_data_log_force[  12] <= 8'h7f;
  filter_in_data_log_force[  13] <= 8'h7f;
  filter_in_data_log_force[  14] <= 8'h7f;
  filter_in_data_log_force[  15] <= 8'h00;
  filter_in_data_log_force[  16] <= 8'h00;
  filter_in_data_log_force[  17] <= 8'h00;
  filter_in_data_log_force[  18] <= 8'h00;
  filter_in_data_log_force[  19] <= 8'h00;
  filter_in_data_log_force[  20] <= 8'h80;
  filter_in_data_log_force[  21] <= 8'h80;
  filter_in_data_log_force[  22] <= 8'h81;
  filter_in_data_log_force[  23] <= 8'h81;
  filter_in_data_log_force[  24] <= 8'h81;
  filter_in_data_log_force[  25] <= 8'h81;
  filter_in_data_log_force[  26] <= 8'h82;
  filter_in_data_log_force[  27] <= 8'h82;
  filter_in_data_log_force[  28] <= 8'h82;
  filter_in_data_log_force[  29] <= 8'h82;
  filter_in_data_log_force[  30] <= 8'h83;
  filter_in_data_log_force[  31] <= 8'h83;
  filter_in_data_log_force[  32] <= 8'h83;
  filter_in_data_log_force[  33] <= 8'h83;
  filter_in_data_log_force[  34] <= 8'h84;
  filter_in_data_log_force[  35] <= 8'h84;
  filter_in_data_log_force[  36] <= 8'h84;
  filter_in_data_log_force[  37] <= 8'h84;
  filter_in_data_log_force[  38] <= 8'h85;
  filter_in_data_log_force[  39] <= 8'h85;
  filter_in_data_log_force[  40] <= 8'h85;
  filter_in_data_log_force[  41] <= 8'h85;
  filter_in_data_log_force[  42] <= 8'h86;
  filter_in_data_log_force[  43] <= 8'h86;
  filter_in_data_log_force[  44] <= 8'h86;
  filter_in_data_log_force[  45] <= 8'h86;
  filter_in_data_log_force[  46] <= 8'h87;
  filter_in_data_log_force[  47] <= 8'h87;
  filter_in_data_log_force[  48] <= 8'h87;
  filter_in_data_log_force[  49] <= 8'h87;
  filter_in_data_log_force[  50] <= 8'h88;
  filter_in_data_log_force[  51] <= 8'h88;
  filter_in_data_log_force[  52] <= 8'h88;
  filter_in_data_log_force[  53] <= 8'h88;
  filter_in_data_log_force[  54] <= 8'h89;
  filter_in_data_log_force[  55] <= 8'h89;
  filter_in_data_log_force[  56] <= 8'h89;
  filter_in_data_log_force[  57] <= 8'h89;
  filter_in_data_log_force[  58] <= 8'h8a;
  filter_in_data_log_force[  59] <= 8'h8a;
  filter_in_data_log_force[  60] <= 8'h8a;
  filter_in_data_log_force[  61] <= 8'h8a;
  filter_in_data_log_force[  62] <= 8'h8b;
  filter_in_data_log_force[  63] <= 8'h8b;
  filter_in_data_log_force[  64] <= 8'h8b;
  filter_in_data_log_force[  65] <= 8'h8b;
  filter_in_data_log_force[  66] <= 8'h8c;
  filter_in_data_log_force[  67] <= 8'h8c;
  filter_in_data_log_force[  68] <= 8'h8c;
  filter_in_data_log_force[  69] <= 8'h8c;
  filter_in_data_log_force[  70] <= 8'h8d;
  filter_in_data_log_force[  71] <= 8'h8d;
  filter_in_data_log_force[  72] <= 8'h8d;
  filter_in_data_log_force[  73] <= 8'h8d;
  filter_in_data_log_force[  74] <= 8'h8e;
  filter_in_data_log_force[  75] <= 8'h8e;
  filter_in_data_log_force[  76] <= 8'h8e;
  filter_in_data_log_force[  77] <= 8'h8e;
  filter_in_data_log_force[  78] <= 8'h8f;
  filter_in_data_log_force[  79] <= 8'h8f;
  filter_in_data_log_force[  80] <= 8'h8f;
  filter_in_data_log_force[  81] <= 8'h8f;
  filter_in_data_log_force[  82] <= 8'h90;
  filter_in_data_log_force[  83] <= 8'h90;
  filter_in_data_log_force[  84] <= 8'h90;
  filter_in_data_log_force[  85] <= 8'h90;
  filter_in_data_log_force[  86] <= 8'h91;
  filter_in_data_log_force[  87] <= 8'h91;
  filter_in_data_log_force[  88] <= 8'h91;
  filter_in_data_log_force[  89] <= 8'h91;
  filter_in_data_log_force[  90] <= 8'h92;
  filter_in_data_log_force[  91] <= 8'h92;
  filter_in_data_log_force[  92] <= 8'h92;
  filter_in_data_log_force[  93] <= 8'h92;
  filter_in_data_log_force[  94] <= 8'h93;
  filter_in_data_log_force[  95] <= 8'h93;
  filter_in_data_log_force[  96] <= 8'h93;
  filter_in_data_log_force[  97] <= 8'h93;
  filter_in_data_log_force[  98] <= 8'h94;
  filter_in_data_log_force[  99] <= 8'h94;
  filter_in_data_log_force[ 100] <= 8'h94;
  filter_in_data_log_force[ 101] <= 8'h94;
  filter_in_data_log_force[ 102] <= 8'h95;
  filter_in_data_log_force[ 103] <= 8'h95;
  filter_in_data_log_force[ 104] <= 8'h95;
  filter_in_data_log_force[ 105] <= 8'h95;
  filter_in_data_log_force[ 106] <= 8'h96;
  filter_in_data_log_force[ 107] <= 8'h96;
  filter_in_data_log_force[ 108] <= 8'h96;
  filter_in_data_log_force[ 109] <= 8'h96;
  filter_in_data_log_force[ 110] <= 8'h97;
  filter_in_data_log_force[ 111] <= 8'h97;
  filter_in_data_log_force[ 112] <= 8'h97;
  filter_in_data_log_force[ 113] <= 8'h97;
  filter_in_data_log_force[ 114] <= 8'h98;
  filter_in_data_log_force[ 115] <= 8'h98;
  filter_in_data_log_force[ 116] <= 8'h98;
  filter_in_data_log_force[ 117] <= 8'h98;
  filter_in_data_log_force[ 118] <= 8'h99;
  filter_in_data_log_force[ 119] <= 8'h99;
  filter_in_data_log_force[ 120] <= 8'h99;
  filter_in_data_log_force[ 121] <= 8'h99;
  filter_in_data_log_force[ 122] <= 8'h9a;
  filter_in_data_log_force[ 123] <= 8'h9a;
  filter_in_data_log_force[ 124] <= 8'h9a;
  filter_in_data_log_force[ 125] <= 8'h9a;
  filter_in_data_log_force[ 126] <= 8'h9b;
  filter_in_data_log_force[ 127] <= 8'h9b;
  filter_in_data_log_force[ 128] <= 8'h9b;
  filter_in_data_log_force[ 129] <= 8'h9b;
  filter_in_data_log_force[ 130] <= 8'h9c;
  filter_in_data_log_force[ 131] <= 8'h9c;
  filter_in_data_log_force[ 132] <= 8'h9c;
  filter_in_data_log_force[ 133] <= 8'h9c;
  filter_in_data_log_force[ 134] <= 8'h9d;
  filter_in_data_log_force[ 135] <= 8'h9d;
  filter_in_data_log_force[ 136] <= 8'h9d;
  filter_in_data_log_force[ 137] <= 8'h9d;
  filter_in_data_log_force[ 138] <= 8'h9e;
  filter_in_data_log_force[ 139] <= 8'h9e;
  filter_in_data_log_force[ 140] <= 8'h9e;
  filter_in_data_log_force[ 141] <= 8'h9e;
  filter_in_data_log_force[ 142] <= 8'h9f;
  filter_in_data_log_force[ 143] <= 8'h9f;
  filter_in_data_log_force[ 144] <= 8'h9f;
  filter_in_data_log_force[ 145] <= 8'h9f;
  filter_in_data_log_force[ 146] <= 8'ha0;
  filter_in_data_log_force[ 147] <= 8'ha0;
  filter_in_data_log_force[ 148] <= 8'ha0;
  filter_in_data_log_force[ 149] <= 8'ha0;
  filter_in_data_log_force[ 150] <= 8'ha1;
  filter_in_data_log_force[ 151] <= 8'ha1;
  filter_in_data_log_force[ 152] <= 8'ha1;
  filter_in_data_log_force[ 153] <= 8'ha1;
  filter_in_data_log_force[ 154] <= 8'ha2;
  filter_in_data_log_force[ 155] <= 8'ha2;
  filter_in_data_log_force[ 156] <= 8'ha2;
  filter_in_data_log_force[ 157] <= 8'ha2;
  filter_in_data_log_force[ 158] <= 8'ha3;
  filter_in_data_log_force[ 159] <= 8'ha3;
  filter_in_data_log_force[ 160] <= 8'ha3;
  filter_in_data_log_force[ 161] <= 8'ha3;
  filter_in_data_log_force[ 162] <= 8'ha4;
  filter_in_data_log_force[ 163] <= 8'ha4;
  filter_in_data_log_force[ 164] <= 8'ha4;
  filter_in_data_log_force[ 165] <= 8'ha4;
  filter_in_data_log_force[ 166] <= 8'ha5;
  filter_in_data_log_force[ 167] <= 8'ha5;
  filter_in_data_log_force[ 168] <= 8'ha5;
  filter_in_data_log_force[ 169] <= 8'ha5;
  filter_in_data_log_force[ 170] <= 8'ha6;
  filter_in_data_log_force[ 171] <= 8'ha6;
  filter_in_data_log_force[ 172] <= 8'ha6;
  filter_in_data_log_force[ 173] <= 8'ha6;
  filter_in_data_log_force[ 174] <= 8'ha7;
  filter_in_data_log_force[ 175] <= 8'ha7;
  filter_in_data_log_force[ 176] <= 8'ha7;
  filter_in_data_log_force[ 177] <= 8'ha7;
  filter_in_data_log_force[ 178] <= 8'ha8;
  filter_in_data_log_force[ 179] <= 8'ha8;
  filter_in_data_log_force[ 180] <= 8'ha8;
  filter_in_data_log_force[ 181] <= 8'ha8;
  filter_in_data_log_force[ 182] <= 8'ha9;
  filter_in_data_log_force[ 183] <= 8'ha9;
  filter_in_data_log_force[ 184] <= 8'ha9;
  filter_in_data_log_force[ 185] <= 8'ha9;
  filter_in_data_log_force[ 186] <= 8'haa;
  filter_in_data_log_force[ 187] <= 8'haa;
  filter_in_data_log_force[ 188] <= 8'haa;
  filter_in_data_log_force[ 189] <= 8'haa;
  filter_in_data_log_force[ 190] <= 8'hab;
  filter_in_data_log_force[ 191] <= 8'hab;
  filter_in_data_log_force[ 192] <= 8'hab;
  filter_in_data_log_force[ 193] <= 8'hab;
  filter_in_data_log_force[ 194] <= 8'hac;
  filter_in_data_log_force[ 195] <= 8'hac;
  filter_in_data_log_force[ 196] <= 8'hac;
  filter_in_data_log_force[ 197] <= 8'hac;
  filter_in_data_log_force[ 198] <= 8'had;
  filter_in_data_log_force[ 199] <= 8'had;
  filter_in_data_log_force[ 200] <= 8'had;
  filter_in_data_log_force[ 201] <= 8'had;
  filter_in_data_log_force[ 202] <= 8'hae;
  filter_in_data_log_force[ 203] <= 8'hae;
  filter_in_data_log_force[ 204] <= 8'hae;
  filter_in_data_log_force[ 205] <= 8'hae;
  filter_in_data_log_force[ 206] <= 8'haf;
  filter_in_data_log_force[ 207] <= 8'haf;
  filter_in_data_log_force[ 208] <= 8'haf;
  filter_in_data_log_force[ 209] <= 8'haf;
  filter_in_data_log_force[ 210] <= 8'hb0;
  filter_in_data_log_force[ 211] <= 8'hb0;
  filter_in_data_log_force[ 212] <= 8'hb0;
  filter_in_data_log_force[ 213] <= 8'hb0;
  filter_in_data_log_force[ 214] <= 8'hb1;
  filter_in_data_log_force[ 215] <= 8'hb1;
  filter_in_data_log_force[ 216] <= 8'hb1;
  filter_in_data_log_force[ 217] <= 8'hb1;
  filter_in_data_log_force[ 218] <= 8'hb2;
  filter_in_data_log_force[ 219] <= 8'hb2;
  filter_in_data_log_force[ 220] <= 8'hb2;
  filter_in_data_log_force[ 221] <= 8'hb2;
  filter_in_data_log_force[ 222] <= 8'hb3;
  filter_in_data_log_force[ 223] <= 8'hb3;
  filter_in_data_log_force[ 224] <= 8'hb3;
  filter_in_data_log_force[ 225] <= 8'hb3;
  filter_in_data_log_force[ 226] <= 8'hb4;
  filter_in_data_log_force[ 227] <= 8'hb4;
  filter_in_data_log_force[ 228] <= 8'hb4;
  filter_in_data_log_force[ 229] <= 8'hb4;
  filter_in_data_log_force[ 230] <= 8'hb5;
  filter_in_data_log_force[ 231] <= 8'hb5;
  filter_in_data_log_force[ 232] <= 8'hb5;
  filter_in_data_log_force[ 233] <= 8'hb5;
  filter_in_data_log_force[ 234] <= 8'hb6;
  filter_in_data_log_force[ 235] <= 8'hb6;
  filter_in_data_log_force[ 236] <= 8'hb6;
  filter_in_data_log_force[ 237] <= 8'hb6;
  filter_in_data_log_force[ 238] <= 8'hb7;
  filter_in_data_log_force[ 239] <= 8'hb7;
  filter_in_data_log_force[ 240] <= 8'hb7;
  filter_in_data_log_force[ 241] <= 8'hb7;
  filter_in_data_log_force[ 242] <= 8'hb8;
  filter_in_data_log_force[ 243] <= 8'hb8;
  filter_in_data_log_force[ 244] <= 8'hb8;
  filter_in_data_log_force[ 245] <= 8'hb8;
  filter_in_data_log_force[ 246] <= 8'hb9;
  filter_in_data_log_force[ 247] <= 8'hb9;
  filter_in_data_log_force[ 248] <= 8'hb9;
  filter_in_data_log_force[ 249] <= 8'hb9;
  filter_in_data_log_force[ 250] <= 8'hba;
  filter_in_data_log_force[ 251] <= 8'hba;
  filter_in_data_log_force[ 252] <= 8'hba;
  filter_in_data_log_force[ 253] <= 8'hba;
  filter_in_data_log_force[ 254] <= 8'hbb;
  filter_in_data_log_force[ 255] <= 8'hbb;
  filter_in_data_log_force[ 256] <= 8'hbb;
  filter_in_data_log_force[ 257] <= 8'hbb;
  filter_in_data_log_force[ 258] <= 8'hbc;
  filter_in_data_log_force[ 259] <= 8'hbc;
  filter_in_data_log_force[ 260] <= 8'hbc;
  filter_in_data_log_force[ 261] <= 8'hbc;
  filter_in_data_log_force[ 262] <= 8'hbd;
  filter_in_data_log_force[ 263] <= 8'hbd;
  filter_in_data_log_force[ 264] <= 8'hbd;
  filter_in_data_log_force[ 265] <= 8'hbd;
  filter_in_data_log_force[ 266] <= 8'hbe;
  filter_in_data_log_force[ 267] <= 8'hbe;
  filter_in_data_log_force[ 268] <= 8'hbe;
  filter_in_data_log_force[ 269] <= 8'hbe;
  filter_in_data_log_force[ 270] <= 8'hbf;
  filter_in_data_log_force[ 271] <= 8'hbf;
  filter_in_data_log_force[ 272] <= 8'hbf;
  filter_in_data_log_force[ 273] <= 8'hbf;
  filter_in_data_log_force[ 274] <= 8'hc0;
  filter_in_data_log_force[ 275] <= 8'hc0;
  filter_in_data_log_force[ 276] <= 8'hc0;
  filter_in_data_log_force[ 277] <= 8'hc0;
  filter_in_data_log_force[ 278] <= 8'hc1;
  filter_in_data_log_force[ 279] <= 8'hc1;
  filter_in_data_log_force[ 280] <= 8'hc1;
  filter_in_data_log_force[ 281] <= 8'hc1;
  filter_in_data_log_force[ 282] <= 8'hc2;
  filter_in_data_log_force[ 283] <= 8'hc2;
  filter_in_data_log_force[ 284] <= 8'hc2;
  filter_in_data_log_force[ 285] <= 8'hc2;
  filter_in_data_log_force[ 286] <= 8'hc3;
  filter_in_data_log_force[ 287] <= 8'hc3;
  filter_in_data_log_force[ 288] <= 8'hc3;
  filter_in_data_log_force[ 289] <= 8'hc3;
  filter_in_data_log_force[ 290] <= 8'hc4;
  filter_in_data_log_force[ 291] <= 8'hc4;
  filter_in_data_log_force[ 292] <= 8'hc4;
  filter_in_data_log_force[ 293] <= 8'hc4;
  filter_in_data_log_force[ 294] <= 8'hc5;
  filter_in_data_log_force[ 295] <= 8'hc5;
  filter_in_data_log_force[ 296] <= 8'hc5;
  filter_in_data_log_force[ 297] <= 8'hc5;
  filter_in_data_log_force[ 298] <= 8'hc6;
  filter_in_data_log_force[ 299] <= 8'hc6;
  filter_in_data_log_force[ 300] <= 8'hc6;
  filter_in_data_log_force[ 301] <= 8'hc6;
  filter_in_data_log_force[ 302] <= 8'hc7;
  filter_in_data_log_force[ 303] <= 8'hc7;
  filter_in_data_log_force[ 304] <= 8'hc7;
  filter_in_data_log_force[ 305] <= 8'hc7;
  filter_in_data_log_force[ 306] <= 8'hc8;
  filter_in_data_log_force[ 307] <= 8'hc8;
  filter_in_data_log_force[ 308] <= 8'hc8;
  filter_in_data_log_force[ 309] <= 8'hc8;
  filter_in_data_log_force[ 310] <= 8'hc9;
  filter_in_data_log_force[ 311] <= 8'hc9;
  filter_in_data_log_force[ 312] <= 8'hc9;
  filter_in_data_log_force[ 313] <= 8'hc9;
  filter_in_data_log_force[ 314] <= 8'hca;
  filter_in_data_log_force[ 315] <= 8'hca;
  filter_in_data_log_force[ 316] <= 8'hca;
  filter_in_data_log_force[ 317] <= 8'hca;
  filter_in_data_log_force[ 318] <= 8'hcb;
  filter_in_data_log_force[ 319] <= 8'hcb;
  filter_in_data_log_force[ 320] <= 8'hcb;
  filter_in_data_log_force[ 321] <= 8'hcb;
  filter_in_data_log_force[ 322] <= 8'hcc;
  filter_in_data_log_force[ 323] <= 8'hcc;
  filter_in_data_log_force[ 324] <= 8'hcc;
  filter_in_data_log_force[ 325] <= 8'hcc;
  filter_in_data_log_force[ 326] <= 8'hcd;
  filter_in_data_log_force[ 327] <= 8'hcd;
  filter_in_data_log_force[ 328] <= 8'hcd;
  filter_in_data_log_force[ 329] <= 8'hcd;
  filter_in_data_log_force[ 330] <= 8'hce;
  filter_in_data_log_force[ 331] <= 8'hce;
  filter_in_data_log_force[ 332] <= 8'hce;
  filter_in_data_log_force[ 333] <= 8'hce;
  filter_in_data_log_force[ 334] <= 8'hcf;
  filter_in_data_log_force[ 335] <= 8'hcf;
  filter_in_data_log_force[ 336] <= 8'hcf;
  filter_in_data_log_force[ 337] <= 8'hcf;
  filter_in_data_log_force[ 338] <= 8'hd0;
  filter_in_data_log_force[ 339] <= 8'hd0;
  filter_in_data_log_force[ 340] <= 8'hd0;
  filter_in_data_log_force[ 341] <= 8'hd0;
  filter_in_data_log_force[ 342] <= 8'hd1;
  filter_in_data_log_force[ 343] <= 8'hd1;
  filter_in_data_log_force[ 344] <= 8'hd1;
  filter_in_data_log_force[ 345] <= 8'hd1;
  filter_in_data_log_force[ 346] <= 8'hd2;
  filter_in_data_log_force[ 347] <= 8'hd2;
  filter_in_data_log_force[ 348] <= 8'hd2;
  filter_in_data_log_force[ 349] <= 8'hd2;
  filter_in_data_log_force[ 350] <= 8'hd3;
  filter_in_data_log_force[ 351] <= 8'hd3;
  filter_in_data_log_force[ 352] <= 8'hd3;
  filter_in_data_log_force[ 353] <= 8'hd3;
  filter_in_data_log_force[ 354] <= 8'hd4;
  filter_in_data_log_force[ 355] <= 8'hd4;
  filter_in_data_log_force[ 356] <= 8'hd4;
  filter_in_data_log_force[ 357] <= 8'hd4;
  filter_in_data_log_force[ 358] <= 8'hd5;
  filter_in_data_log_force[ 359] <= 8'hd5;
  filter_in_data_log_force[ 360] <= 8'hd5;
  filter_in_data_log_force[ 361] <= 8'hd5;
  filter_in_data_log_force[ 362] <= 8'hd6;
  filter_in_data_log_force[ 363] <= 8'hd6;
  filter_in_data_log_force[ 364] <= 8'hd6;
  filter_in_data_log_force[ 365] <= 8'hd6;
  filter_in_data_log_force[ 366] <= 8'hd7;
  filter_in_data_log_force[ 367] <= 8'hd7;
  filter_in_data_log_force[ 368] <= 8'hd7;
  filter_in_data_log_force[ 369] <= 8'hd7;
  filter_in_data_log_force[ 370] <= 8'hd8;
  filter_in_data_log_force[ 371] <= 8'hd8;
  filter_in_data_log_force[ 372] <= 8'hd8;
  filter_in_data_log_force[ 373] <= 8'hd8;
  filter_in_data_log_force[ 374] <= 8'hd9;
  filter_in_data_log_force[ 375] <= 8'hd9;
  filter_in_data_log_force[ 376] <= 8'hd9;
  filter_in_data_log_force[ 377] <= 8'hd9;
  filter_in_data_log_force[ 378] <= 8'hda;
  filter_in_data_log_force[ 379] <= 8'hda;
  filter_in_data_log_force[ 380] <= 8'hda;
  filter_in_data_log_force[ 381] <= 8'hda;
  filter_in_data_log_force[ 382] <= 8'hdb;
  filter_in_data_log_force[ 383] <= 8'hdb;
  filter_in_data_log_force[ 384] <= 8'hdb;
  filter_in_data_log_force[ 385] <= 8'hdb;
  filter_in_data_log_force[ 386] <= 8'hdc;
  filter_in_data_log_force[ 387] <= 8'hdc;
  filter_in_data_log_force[ 388] <= 8'hdc;
  filter_in_data_log_force[ 389] <= 8'hdc;
  filter_in_data_log_force[ 390] <= 8'hdd;
  filter_in_data_log_force[ 391] <= 8'hdd;
  filter_in_data_log_force[ 392] <= 8'hdd;
  filter_in_data_log_force[ 393] <= 8'hdd;
  filter_in_data_log_force[ 394] <= 8'hde;
  filter_in_data_log_force[ 395] <= 8'hde;
  filter_in_data_log_force[ 396] <= 8'hde;
  filter_in_data_log_force[ 397] <= 8'hde;
  filter_in_data_log_force[ 398] <= 8'hdf;
  filter_in_data_log_force[ 399] <= 8'hdf;
  filter_in_data_log_force[ 400] <= 8'hdf;
  filter_in_data_log_force[ 401] <= 8'hdf;
  filter_in_data_log_force[ 402] <= 8'he0;
  filter_in_data_log_force[ 403] <= 8'he0;
  filter_in_data_log_force[ 404] <= 8'he0;
  filter_in_data_log_force[ 405] <= 8'he0;
  filter_in_data_log_force[ 406] <= 8'he1;
  filter_in_data_log_force[ 407] <= 8'he1;
  filter_in_data_log_force[ 408] <= 8'he1;
  filter_in_data_log_force[ 409] <= 8'he1;
  filter_in_data_log_force[ 410] <= 8'he2;
  filter_in_data_log_force[ 411] <= 8'he2;
  filter_in_data_log_force[ 412] <= 8'he2;
  filter_in_data_log_force[ 413] <= 8'he2;
  filter_in_data_log_force[ 414] <= 8'he3;
  filter_in_data_log_force[ 415] <= 8'he3;
  filter_in_data_log_force[ 416] <= 8'he3;
  filter_in_data_log_force[ 417] <= 8'he3;
  filter_in_data_log_force[ 418] <= 8'he4;
  filter_in_data_log_force[ 419] <= 8'he4;
  filter_in_data_log_force[ 420] <= 8'he4;
  filter_in_data_log_force[ 421] <= 8'he4;
  filter_in_data_log_force[ 422] <= 8'he5;
  filter_in_data_log_force[ 423] <= 8'he5;
  filter_in_data_log_force[ 424] <= 8'he5;
  filter_in_data_log_force[ 425] <= 8'he5;
  filter_in_data_log_force[ 426] <= 8'he6;
  filter_in_data_log_force[ 427] <= 8'he6;
  filter_in_data_log_force[ 428] <= 8'he6;
  filter_in_data_log_force[ 429] <= 8'he6;
  filter_in_data_log_force[ 430] <= 8'he7;
  filter_in_data_log_force[ 431] <= 8'he7;
  filter_in_data_log_force[ 432] <= 8'he7;
  filter_in_data_log_force[ 433] <= 8'he7;
  filter_in_data_log_force[ 434] <= 8'he8;
  filter_in_data_log_force[ 435] <= 8'he8;
  filter_in_data_log_force[ 436] <= 8'he8;
  filter_in_data_log_force[ 437] <= 8'he8;
  filter_in_data_log_force[ 438] <= 8'he9;
  filter_in_data_log_force[ 439] <= 8'he9;
  filter_in_data_log_force[ 440] <= 8'he9;
  filter_in_data_log_force[ 441] <= 8'he9;
  filter_in_data_log_force[ 442] <= 8'hea;
  filter_in_data_log_force[ 443] <= 8'hea;
  filter_in_data_log_force[ 444] <= 8'hea;
  filter_in_data_log_force[ 445] <= 8'hea;
  filter_in_data_log_force[ 446] <= 8'heb;
  filter_in_data_log_force[ 447] <= 8'heb;
  filter_in_data_log_force[ 448] <= 8'heb;
  filter_in_data_log_force[ 449] <= 8'heb;
  filter_in_data_log_force[ 450] <= 8'hec;
  filter_in_data_log_force[ 451] <= 8'hec;
  filter_in_data_log_force[ 452] <= 8'hec;
  filter_in_data_log_force[ 453] <= 8'hec;
  filter_in_data_log_force[ 454] <= 8'hed;
  filter_in_data_log_force[ 455] <= 8'hed;
  filter_in_data_log_force[ 456] <= 8'hed;
  filter_in_data_log_force[ 457] <= 8'hed;
  filter_in_data_log_force[ 458] <= 8'hee;
  filter_in_data_log_force[ 459] <= 8'hee;
  filter_in_data_log_force[ 460] <= 8'hee;
  filter_in_data_log_force[ 461] <= 8'hee;
  filter_in_data_log_force[ 462] <= 8'hef;
  filter_in_data_log_force[ 463] <= 8'hef;
  filter_in_data_log_force[ 464] <= 8'hef;
  filter_in_data_log_force[ 465] <= 8'hef;
  filter_in_data_log_force[ 466] <= 8'hf0;
  filter_in_data_log_force[ 467] <= 8'hf0;
  filter_in_data_log_force[ 468] <= 8'hf0;
  filter_in_data_log_force[ 469] <= 8'hf0;
  filter_in_data_log_force[ 470] <= 8'hf1;
  filter_in_data_log_force[ 471] <= 8'hf1;
  filter_in_data_log_force[ 472] <= 8'hf1;
  filter_in_data_log_force[ 473] <= 8'hf1;
  filter_in_data_log_force[ 474] <= 8'hf2;
  filter_in_data_log_force[ 475] <= 8'hf2;
  filter_in_data_log_force[ 476] <= 8'hf2;
  filter_in_data_log_force[ 477] <= 8'hf2;
  filter_in_data_log_force[ 478] <= 8'hf3;
  filter_in_data_log_force[ 479] <= 8'hf3;
  filter_in_data_log_force[ 480] <= 8'hf3;
  filter_in_data_log_force[ 481] <= 8'hf3;
  filter_in_data_log_force[ 482] <= 8'hf4;
  filter_in_data_log_force[ 483] <= 8'hf4;
  filter_in_data_log_force[ 484] <= 8'hf4;
  filter_in_data_log_force[ 485] <= 8'hf4;
  filter_in_data_log_force[ 486] <= 8'hf5;
  filter_in_data_log_force[ 487] <= 8'hf5;
  filter_in_data_log_force[ 488] <= 8'hf5;
  filter_in_data_log_force[ 489] <= 8'hf5;
  filter_in_data_log_force[ 490] <= 8'hf6;
  filter_in_data_log_force[ 491] <= 8'hf6;
  filter_in_data_log_force[ 492] <= 8'hf6;
  filter_in_data_log_force[ 493] <= 8'hf6;
  filter_in_data_log_force[ 494] <= 8'hf7;
  filter_in_data_log_force[ 495] <= 8'hf7;
  filter_in_data_log_force[ 496] <= 8'hf7;
  filter_in_data_log_force[ 497] <= 8'hf7;
  filter_in_data_log_force[ 498] <= 8'hf8;
  filter_in_data_log_force[ 499] <= 8'hf8;
  filter_in_data_log_force[ 500] <= 8'hf8;
  filter_in_data_log_force[ 501] <= 8'hf8;
  filter_in_data_log_force[ 502] <= 8'hf9;
  filter_in_data_log_force[ 503] <= 8'hf9;
  filter_in_data_log_force[ 504] <= 8'hf9;
  filter_in_data_log_force[ 505] <= 8'hf9;
  filter_in_data_log_force[ 506] <= 8'hfa;
  filter_in_data_log_force[ 507] <= 8'hfa;
  filter_in_data_log_force[ 508] <= 8'hfa;
  filter_in_data_log_force[ 509] <= 8'hfa;
  filter_in_data_log_force[ 510] <= 8'hfb;
  filter_in_data_log_force[ 511] <= 8'hfb;
  filter_in_data_log_force[ 512] <= 8'hfb;
  filter_in_data_log_force[ 513] <= 8'hfb;
  filter_in_data_log_force[ 514] <= 8'hfc;
  filter_in_data_log_force[ 515] <= 8'hfc;
  filter_in_data_log_force[ 516] <= 8'hfc;
  filter_in_data_log_force[ 517] <= 8'hfc;
  filter_in_data_log_force[ 518] <= 8'hfd;
  filter_in_data_log_force[ 519] <= 8'hfd;
  filter_in_data_log_force[ 520] <= 8'hfd;
  filter_in_data_log_force[ 521] <= 8'hfd;
  filter_in_data_log_force[ 522] <= 8'hfe;
  filter_in_data_log_force[ 523] <= 8'hfe;
  filter_in_data_log_force[ 524] <= 8'hfe;
  filter_in_data_log_force[ 525] <= 8'hfe;
  filter_in_data_log_force[ 526] <= 8'hff;
  filter_in_data_log_force[ 527] <= 8'hff;
  filter_in_data_log_force[ 528] <= 8'hff;
  filter_in_data_log_force[ 529] <= 8'hff;
  filter_in_data_log_force[ 530] <= 8'h00;
  filter_in_data_log_force[ 531] <= 8'h00;
  filter_in_data_log_force[ 532] <= 8'h00;
  filter_in_data_log_force[ 533] <= 8'h00;
  filter_in_data_log_force[ 534] <= 8'h01;
  filter_in_data_log_force[ 535] <= 8'h01;
  filter_in_data_log_force[ 536] <= 8'h01;
  filter_in_data_log_force[ 537] <= 8'h01;
  filter_in_data_log_force[ 538] <= 8'h02;
  filter_in_data_log_force[ 539] <= 8'h02;
  filter_in_data_log_force[ 540] <= 8'h02;
  filter_in_data_log_force[ 541] <= 8'h02;
  filter_in_data_log_force[ 542] <= 8'h03;
  filter_in_data_log_force[ 543] <= 8'h03;
  filter_in_data_log_force[ 544] <= 8'h03;
  filter_in_data_log_force[ 545] <= 8'h03;
  filter_in_data_log_force[ 546] <= 8'h04;
  filter_in_data_log_force[ 547] <= 8'h04;
  filter_in_data_log_force[ 548] <= 8'h04;
  filter_in_data_log_force[ 549] <= 8'h04;
  filter_in_data_log_force[ 550] <= 8'h05;
  filter_in_data_log_force[ 551] <= 8'h05;
  filter_in_data_log_force[ 552] <= 8'h05;
  filter_in_data_log_force[ 553] <= 8'h05;
  filter_in_data_log_force[ 554] <= 8'h06;
  filter_in_data_log_force[ 555] <= 8'h06;
  filter_in_data_log_force[ 556] <= 8'h06;
  filter_in_data_log_force[ 557] <= 8'h06;
  filter_in_data_log_force[ 558] <= 8'h07;
  filter_in_data_log_force[ 559] <= 8'h07;
  filter_in_data_log_force[ 560] <= 8'h07;
  filter_in_data_log_force[ 561] <= 8'h07;
  filter_in_data_log_force[ 562] <= 8'h08;
  filter_in_data_log_force[ 563] <= 8'h08;
  filter_in_data_log_force[ 564] <= 8'h08;
  filter_in_data_log_force[ 565] <= 8'h08;
  filter_in_data_log_force[ 566] <= 8'h09;
  filter_in_data_log_force[ 567] <= 8'h09;
  filter_in_data_log_force[ 568] <= 8'h09;
  filter_in_data_log_force[ 569] <= 8'h09;
  filter_in_data_log_force[ 570] <= 8'h0a;
  filter_in_data_log_force[ 571] <= 8'h0a;
  filter_in_data_log_force[ 572] <= 8'h0a;
  filter_in_data_log_force[ 573] <= 8'h0a;
  filter_in_data_log_force[ 574] <= 8'h0b;
  filter_in_data_log_force[ 575] <= 8'h0b;
  filter_in_data_log_force[ 576] <= 8'h0b;
  filter_in_data_log_force[ 577] <= 8'h0b;
  filter_in_data_log_force[ 578] <= 8'h0c;
  filter_in_data_log_force[ 579] <= 8'h0c;
  filter_in_data_log_force[ 580] <= 8'h0c;
  filter_in_data_log_force[ 581] <= 8'h0c;
  filter_in_data_log_force[ 582] <= 8'h0d;
  filter_in_data_log_force[ 583] <= 8'h0d;
  filter_in_data_log_force[ 584] <= 8'h0d;
  filter_in_data_log_force[ 585] <= 8'h0d;
  filter_in_data_log_force[ 586] <= 8'h0e;
  filter_in_data_log_force[ 587] <= 8'h0e;
  filter_in_data_log_force[ 588] <= 8'h0e;
  filter_in_data_log_force[ 589] <= 8'h0e;
  filter_in_data_log_force[ 590] <= 8'h0f;
  filter_in_data_log_force[ 591] <= 8'h0f;
  filter_in_data_log_force[ 592] <= 8'h0f;
  filter_in_data_log_force[ 593] <= 8'h0f;
  filter_in_data_log_force[ 594] <= 8'h10;
  filter_in_data_log_force[ 595] <= 8'h10;
  filter_in_data_log_force[ 596] <= 8'h10;
  filter_in_data_log_force[ 597] <= 8'h10;
  filter_in_data_log_force[ 598] <= 8'h11;
  filter_in_data_log_force[ 599] <= 8'h11;
  filter_in_data_log_force[ 600] <= 8'h11;
  filter_in_data_log_force[ 601] <= 8'h11;
  filter_in_data_log_force[ 602] <= 8'h12;
  filter_in_data_log_force[ 603] <= 8'h12;
  filter_in_data_log_force[ 604] <= 8'h12;
  filter_in_data_log_force[ 605] <= 8'h12;
  filter_in_data_log_force[ 606] <= 8'h13;
  filter_in_data_log_force[ 607] <= 8'h13;
  filter_in_data_log_force[ 608] <= 8'h13;
  filter_in_data_log_force[ 609] <= 8'h13;
  filter_in_data_log_force[ 610] <= 8'h14;
  filter_in_data_log_force[ 611] <= 8'h14;
  filter_in_data_log_force[ 612] <= 8'h14;
  filter_in_data_log_force[ 613] <= 8'h14;
  filter_in_data_log_force[ 614] <= 8'h15;
  filter_in_data_log_force[ 615] <= 8'h15;
  filter_in_data_log_force[ 616] <= 8'h15;
  filter_in_data_log_force[ 617] <= 8'h15;
  filter_in_data_log_force[ 618] <= 8'h16;
  filter_in_data_log_force[ 619] <= 8'h16;
  filter_in_data_log_force[ 620] <= 8'h16;
  filter_in_data_log_force[ 621] <= 8'h16;
  filter_in_data_log_force[ 622] <= 8'h17;
  filter_in_data_log_force[ 623] <= 8'h17;
  filter_in_data_log_force[ 624] <= 8'h17;
  filter_in_data_log_force[ 625] <= 8'h17;
  filter_in_data_log_force[ 626] <= 8'h18;
  filter_in_data_log_force[ 627] <= 8'h18;
  filter_in_data_log_force[ 628] <= 8'h18;
  filter_in_data_log_force[ 629] <= 8'h18;
  filter_in_data_log_force[ 630] <= 8'h19;
  filter_in_data_log_force[ 631] <= 8'h19;
  filter_in_data_log_force[ 632] <= 8'h19;
  filter_in_data_log_force[ 633] <= 8'h19;
  filter_in_data_log_force[ 634] <= 8'h1a;
  filter_in_data_log_force[ 635] <= 8'h1a;
  filter_in_data_log_force[ 636] <= 8'h1a;
  filter_in_data_log_force[ 637] <= 8'h1a;
  filter_in_data_log_force[ 638] <= 8'h1b;
  filter_in_data_log_force[ 639] <= 8'h1b;
  filter_in_data_log_force[ 640] <= 8'h1b;
  filter_in_data_log_force[ 641] <= 8'h1b;
  filter_in_data_log_force[ 642] <= 8'h1c;
  filter_in_data_log_force[ 643] <= 8'h1c;
  filter_in_data_log_force[ 644] <= 8'h1c;
  filter_in_data_log_force[ 645] <= 8'h1c;
  filter_in_data_log_force[ 646] <= 8'h1d;
  filter_in_data_log_force[ 647] <= 8'h1d;
  filter_in_data_log_force[ 648] <= 8'h1d;
  filter_in_data_log_force[ 649] <= 8'h1d;
  filter_in_data_log_force[ 650] <= 8'h1e;
  filter_in_data_log_force[ 651] <= 8'h1e;
  filter_in_data_log_force[ 652] <= 8'h1e;
  filter_in_data_log_force[ 653] <= 8'h1e;
  filter_in_data_log_force[ 654] <= 8'h1f;
  filter_in_data_log_force[ 655] <= 8'h1f;
  filter_in_data_log_force[ 656] <= 8'h1f;
  filter_in_data_log_force[ 657] <= 8'h1f;
  filter_in_data_log_force[ 658] <= 8'h20;
  filter_in_data_log_force[ 659] <= 8'h20;
  filter_in_data_log_force[ 660] <= 8'h20;
  filter_in_data_log_force[ 661] <= 8'h20;
  filter_in_data_log_force[ 662] <= 8'h21;
  filter_in_data_log_force[ 663] <= 8'h21;
  filter_in_data_log_force[ 664] <= 8'h21;
  filter_in_data_log_force[ 665] <= 8'h21;
  filter_in_data_log_force[ 666] <= 8'h22;
  filter_in_data_log_force[ 667] <= 8'h22;
  filter_in_data_log_force[ 668] <= 8'h22;
  filter_in_data_log_force[ 669] <= 8'h22;
  filter_in_data_log_force[ 670] <= 8'h23;
  filter_in_data_log_force[ 671] <= 8'h23;
  filter_in_data_log_force[ 672] <= 8'h23;
  filter_in_data_log_force[ 673] <= 8'h23;
  filter_in_data_log_force[ 674] <= 8'h24;
  filter_in_data_log_force[ 675] <= 8'h24;
  filter_in_data_log_force[ 676] <= 8'h24;
  filter_in_data_log_force[ 677] <= 8'h24;
  filter_in_data_log_force[ 678] <= 8'h25;
  filter_in_data_log_force[ 679] <= 8'h25;
  filter_in_data_log_force[ 680] <= 8'h25;
  filter_in_data_log_force[ 681] <= 8'h25;
  filter_in_data_log_force[ 682] <= 8'h26;
  filter_in_data_log_force[ 683] <= 8'h26;
  filter_in_data_log_force[ 684] <= 8'h26;
  filter_in_data_log_force[ 685] <= 8'h26;
  filter_in_data_log_force[ 686] <= 8'h27;
  filter_in_data_log_force[ 687] <= 8'h27;
  filter_in_data_log_force[ 688] <= 8'h27;
  filter_in_data_log_force[ 689] <= 8'h27;
  filter_in_data_log_force[ 690] <= 8'h28;
  filter_in_data_log_force[ 691] <= 8'h28;
  filter_in_data_log_force[ 692] <= 8'h28;
  filter_in_data_log_force[ 693] <= 8'h28;
  filter_in_data_log_force[ 694] <= 8'h29;
  filter_in_data_log_force[ 695] <= 8'h29;
  filter_in_data_log_force[ 696] <= 8'h29;
  filter_in_data_log_force[ 697] <= 8'h29;
  filter_in_data_log_force[ 698] <= 8'h2a;
  filter_in_data_log_force[ 699] <= 8'h2a;
  filter_in_data_log_force[ 700] <= 8'h2a;
  filter_in_data_log_force[ 701] <= 8'h2a;
  filter_in_data_log_force[ 702] <= 8'h2b;
  filter_in_data_log_force[ 703] <= 8'h2b;
  filter_in_data_log_force[ 704] <= 8'h2b;
  filter_in_data_log_force[ 705] <= 8'h2b;
  filter_in_data_log_force[ 706] <= 8'h2c;
  filter_in_data_log_force[ 707] <= 8'h2c;
  filter_in_data_log_force[ 708] <= 8'h2c;
  filter_in_data_log_force[ 709] <= 8'h2c;
  filter_in_data_log_force[ 710] <= 8'h2d;
  filter_in_data_log_force[ 711] <= 8'h2d;
  filter_in_data_log_force[ 712] <= 8'h2d;
  filter_in_data_log_force[ 713] <= 8'h2d;
  filter_in_data_log_force[ 714] <= 8'h2e;
  filter_in_data_log_force[ 715] <= 8'h2e;
  filter_in_data_log_force[ 716] <= 8'h2e;
  filter_in_data_log_force[ 717] <= 8'h2e;
  filter_in_data_log_force[ 718] <= 8'h2f;
  filter_in_data_log_force[ 719] <= 8'h2f;
  filter_in_data_log_force[ 720] <= 8'h2f;
  filter_in_data_log_force[ 721] <= 8'h2f;
  filter_in_data_log_force[ 722] <= 8'h30;
  filter_in_data_log_force[ 723] <= 8'h30;
  filter_in_data_log_force[ 724] <= 8'h30;
  filter_in_data_log_force[ 725] <= 8'h30;
  filter_in_data_log_force[ 726] <= 8'h31;
  filter_in_data_log_force[ 727] <= 8'h31;
  filter_in_data_log_force[ 728] <= 8'h31;
  filter_in_data_log_force[ 729] <= 8'h31;
  filter_in_data_log_force[ 730] <= 8'h32;
  filter_in_data_log_force[ 731] <= 8'h32;
  filter_in_data_log_force[ 732] <= 8'h32;
  filter_in_data_log_force[ 733] <= 8'h32;
  filter_in_data_log_force[ 734] <= 8'h33;
  filter_in_data_log_force[ 735] <= 8'h33;
  filter_in_data_log_force[ 736] <= 8'h33;
  filter_in_data_log_force[ 737] <= 8'h33;
  filter_in_data_log_force[ 738] <= 8'h34;
  filter_in_data_log_force[ 739] <= 8'h34;
  filter_in_data_log_force[ 740] <= 8'h34;
  filter_in_data_log_force[ 741] <= 8'h34;
  filter_in_data_log_force[ 742] <= 8'h35;
  filter_in_data_log_force[ 743] <= 8'h35;
  filter_in_data_log_force[ 744] <= 8'h35;
  filter_in_data_log_force[ 745] <= 8'h35;
  filter_in_data_log_force[ 746] <= 8'h36;
  filter_in_data_log_force[ 747] <= 8'h36;
  filter_in_data_log_force[ 748] <= 8'h36;
  filter_in_data_log_force[ 749] <= 8'h36;
  filter_in_data_log_force[ 750] <= 8'h37;
  filter_in_data_log_force[ 751] <= 8'h37;
  filter_in_data_log_force[ 752] <= 8'h37;
  filter_in_data_log_force[ 753] <= 8'h37;
  filter_in_data_log_force[ 754] <= 8'h38;
  filter_in_data_log_force[ 755] <= 8'h38;
  filter_in_data_log_force[ 756] <= 8'h38;
  filter_in_data_log_force[ 757] <= 8'h38;
  filter_in_data_log_force[ 758] <= 8'h39;
  filter_in_data_log_force[ 759] <= 8'h39;
  filter_in_data_log_force[ 760] <= 8'h39;
  filter_in_data_log_force[ 761] <= 8'h39;
  filter_in_data_log_force[ 762] <= 8'h3a;
  filter_in_data_log_force[ 763] <= 8'h3a;
  filter_in_data_log_force[ 764] <= 8'h3a;
  filter_in_data_log_force[ 765] <= 8'h3a;
  filter_in_data_log_force[ 766] <= 8'h3b;
  filter_in_data_log_force[ 767] <= 8'h3b;
  filter_in_data_log_force[ 768] <= 8'h3b;
  filter_in_data_log_force[ 769] <= 8'h3b;
  filter_in_data_log_force[ 770] <= 8'h3c;
  filter_in_data_log_force[ 771] <= 8'h3c;
  filter_in_data_log_force[ 772] <= 8'h3c;
  filter_in_data_log_force[ 773] <= 8'h3c;
  filter_in_data_log_force[ 774] <= 8'h3d;
  filter_in_data_log_force[ 775] <= 8'h3d;
  filter_in_data_log_force[ 776] <= 8'h3d;
  filter_in_data_log_force[ 777] <= 8'h3d;
  filter_in_data_log_force[ 778] <= 8'h3e;
  filter_in_data_log_force[ 779] <= 8'h3e;
  filter_in_data_log_force[ 780] <= 8'h3e;
  filter_in_data_log_force[ 781] <= 8'h3e;
  filter_in_data_log_force[ 782] <= 8'h3f;
  filter_in_data_log_force[ 783] <= 8'h3f;
  filter_in_data_log_force[ 784] <= 8'h3f;
  filter_in_data_log_force[ 785] <= 8'h3f;
  filter_in_data_log_force[ 786] <= 8'h40;
  filter_in_data_log_force[ 787] <= 8'h40;
  filter_in_data_log_force[ 788] <= 8'h40;
  filter_in_data_log_force[ 789] <= 8'h40;
  filter_in_data_log_force[ 790] <= 8'h41;
  filter_in_data_log_force[ 791] <= 8'h41;
  filter_in_data_log_force[ 792] <= 8'h41;
  filter_in_data_log_force[ 793] <= 8'h41;
  filter_in_data_log_force[ 794] <= 8'h42;
  filter_in_data_log_force[ 795] <= 8'h42;
  filter_in_data_log_force[ 796] <= 8'h42;
  filter_in_data_log_force[ 797] <= 8'h42;
  filter_in_data_log_force[ 798] <= 8'h43;
  filter_in_data_log_force[ 799] <= 8'h43;
  filter_in_data_log_force[ 800] <= 8'h43;
  filter_in_data_log_force[ 801] <= 8'h43;
  filter_in_data_log_force[ 802] <= 8'h44;
  filter_in_data_log_force[ 803] <= 8'h44;
  filter_in_data_log_force[ 804] <= 8'h44;
  filter_in_data_log_force[ 805] <= 8'h44;
  filter_in_data_log_force[ 806] <= 8'h45;
  filter_in_data_log_force[ 807] <= 8'h45;
  filter_in_data_log_force[ 808] <= 8'h45;
  filter_in_data_log_force[ 809] <= 8'h45;
  filter_in_data_log_force[ 810] <= 8'h46;
  filter_in_data_log_force[ 811] <= 8'h46;
  filter_in_data_log_force[ 812] <= 8'h46;
  filter_in_data_log_force[ 813] <= 8'h46;
  filter_in_data_log_force[ 814] <= 8'h47;
  filter_in_data_log_force[ 815] <= 8'h47;
  filter_in_data_log_force[ 816] <= 8'h47;
  filter_in_data_log_force[ 817] <= 8'h47;
  filter_in_data_log_force[ 818] <= 8'h48;
  filter_in_data_log_force[ 819] <= 8'h48;
  filter_in_data_log_force[ 820] <= 8'h48;
  filter_in_data_log_force[ 821] <= 8'h48;
  filter_in_data_log_force[ 822] <= 8'h49;
  filter_in_data_log_force[ 823] <= 8'h49;
  filter_in_data_log_force[ 824] <= 8'h49;
  filter_in_data_log_force[ 825] <= 8'h49;
  filter_in_data_log_force[ 826] <= 8'h4a;
  filter_in_data_log_force[ 827] <= 8'h4a;
  filter_in_data_log_force[ 828] <= 8'h4a;
  filter_in_data_log_force[ 829] <= 8'h4a;
  filter_in_data_log_force[ 830] <= 8'h4b;
  filter_in_data_log_force[ 831] <= 8'h4b;
  filter_in_data_log_force[ 832] <= 8'h4b;
  filter_in_data_log_force[ 833] <= 8'h4b;
  filter_in_data_log_force[ 834] <= 8'h4c;
  filter_in_data_log_force[ 835] <= 8'h4c;
  filter_in_data_log_force[ 836] <= 8'h4c;
  filter_in_data_log_force[ 837] <= 8'h4c;
  filter_in_data_log_force[ 838] <= 8'h4d;
  filter_in_data_log_force[ 839] <= 8'h4d;
  filter_in_data_log_force[ 840] <= 8'h4d;
  filter_in_data_log_force[ 841] <= 8'h4d;
  filter_in_data_log_force[ 842] <= 8'h4e;
  filter_in_data_log_force[ 843] <= 8'h4e;
  filter_in_data_log_force[ 844] <= 8'h4e;
  filter_in_data_log_force[ 845] <= 8'h4e;
  filter_in_data_log_force[ 846] <= 8'h4f;
  filter_in_data_log_force[ 847] <= 8'h4f;
  filter_in_data_log_force[ 848] <= 8'h4f;
  filter_in_data_log_force[ 849] <= 8'h4f;
  filter_in_data_log_force[ 850] <= 8'h50;
  filter_in_data_log_force[ 851] <= 8'h50;
  filter_in_data_log_force[ 852] <= 8'h50;
  filter_in_data_log_force[ 853] <= 8'h50;
  filter_in_data_log_force[ 854] <= 8'h51;
  filter_in_data_log_force[ 855] <= 8'h51;
  filter_in_data_log_force[ 856] <= 8'h51;
  filter_in_data_log_force[ 857] <= 8'h51;
  filter_in_data_log_force[ 858] <= 8'h52;
  filter_in_data_log_force[ 859] <= 8'h52;
  filter_in_data_log_force[ 860] <= 8'h52;
  filter_in_data_log_force[ 861] <= 8'h52;
  filter_in_data_log_force[ 862] <= 8'h53;
  filter_in_data_log_force[ 863] <= 8'h53;
  filter_in_data_log_force[ 864] <= 8'h53;
  filter_in_data_log_force[ 865] <= 8'h53;
  filter_in_data_log_force[ 866] <= 8'h54;
  filter_in_data_log_force[ 867] <= 8'h54;
  filter_in_data_log_force[ 868] <= 8'h54;
  filter_in_data_log_force[ 869] <= 8'h54;
  filter_in_data_log_force[ 870] <= 8'h55;
  filter_in_data_log_force[ 871] <= 8'h55;
  filter_in_data_log_force[ 872] <= 8'h55;
  filter_in_data_log_force[ 873] <= 8'h55;
  filter_in_data_log_force[ 874] <= 8'h56;
  filter_in_data_log_force[ 875] <= 8'h56;
  filter_in_data_log_force[ 876] <= 8'h56;
  filter_in_data_log_force[ 877] <= 8'h56;
  filter_in_data_log_force[ 878] <= 8'h57;
  filter_in_data_log_force[ 879] <= 8'h57;
  filter_in_data_log_force[ 880] <= 8'h57;
  filter_in_data_log_force[ 881] <= 8'h57;
  filter_in_data_log_force[ 882] <= 8'h58;
  filter_in_data_log_force[ 883] <= 8'h58;
  filter_in_data_log_force[ 884] <= 8'h58;
  filter_in_data_log_force[ 885] <= 8'h58;
  filter_in_data_log_force[ 886] <= 8'h59;
  filter_in_data_log_force[ 887] <= 8'h59;
  filter_in_data_log_force[ 888] <= 8'h59;
  filter_in_data_log_force[ 889] <= 8'h59;
  filter_in_data_log_force[ 890] <= 8'h5a;
  filter_in_data_log_force[ 891] <= 8'h5a;
  filter_in_data_log_force[ 892] <= 8'h5a;
  filter_in_data_log_force[ 893] <= 8'h5a;
  filter_in_data_log_force[ 894] <= 8'h5b;
  filter_in_data_log_force[ 895] <= 8'h5b;
  filter_in_data_log_force[ 896] <= 8'h5b;
  filter_in_data_log_force[ 897] <= 8'h5b;
  filter_in_data_log_force[ 898] <= 8'h5c;
  filter_in_data_log_force[ 899] <= 8'h5c;
  filter_in_data_log_force[ 900] <= 8'h5c;
  filter_in_data_log_force[ 901] <= 8'h5c;
  filter_in_data_log_force[ 902] <= 8'h5d;
  filter_in_data_log_force[ 903] <= 8'h5d;
  filter_in_data_log_force[ 904] <= 8'h5d;
  filter_in_data_log_force[ 905] <= 8'h5d;
  filter_in_data_log_force[ 906] <= 8'h5e;
  filter_in_data_log_force[ 907] <= 8'h5e;
  filter_in_data_log_force[ 908] <= 8'h5e;
  filter_in_data_log_force[ 909] <= 8'h5e;
  filter_in_data_log_force[ 910] <= 8'h5f;
  filter_in_data_log_force[ 911] <= 8'h5f;
  filter_in_data_log_force[ 912] <= 8'h5f;
  filter_in_data_log_force[ 913] <= 8'h5f;
  filter_in_data_log_force[ 914] <= 8'h60;
  filter_in_data_log_force[ 915] <= 8'h60;
  filter_in_data_log_force[ 916] <= 8'h60;
  filter_in_data_log_force[ 917] <= 8'h60;
  filter_in_data_log_force[ 918] <= 8'h61;
  filter_in_data_log_force[ 919] <= 8'h61;
  filter_in_data_log_force[ 920] <= 8'h61;
  filter_in_data_log_force[ 921] <= 8'h61;
  filter_in_data_log_force[ 922] <= 8'h62;
  filter_in_data_log_force[ 923] <= 8'h62;
  filter_in_data_log_force[ 924] <= 8'h62;
  filter_in_data_log_force[ 925] <= 8'h62;
  filter_in_data_log_force[ 926] <= 8'h63;
  filter_in_data_log_force[ 927] <= 8'h63;
  filter_in_data_log_force[ 928] <= 8'h63;
  filter_in_data_log_force[ 929] <= 8'h63;
  filter_in_data_log_force[ 930] <= 8'h64;
  filter_in_data_log_force[ 931] <= 8'h64;
  filter_in_data_log_force[ 932] <= 8'h64;
  filter_in_data_log_force[ 933] <= 8'h64;
  filter_in_data_log_force[ 934] <= 8'h65;
  filter_in_data_log_force[ 935] <= 8'h65;
  filter_in_data_log_force[ 936] <= 8'h65;
  filter_in_data_log_force[ 937] <= 8'h65;
  filter_in_data_log_force[ 938] <= 8'h66;
  filter_in_data_log_force[ 939] <= 8'h66;
  filter_in_data_log_force[ 940] <= 8'h66;
  filter_in_data_log_force[ 941] <= 8'h66;
  filter_in_data_log_force[ 942] <= 8'h67;
  filter_in_data_log_force[ 943] <= 8'h67;
  filter_in_data_log_force[ 944] <= 8'h67;
  filter_in_data_log_force[ 945] <= 8'h67;
  filter_in_data_log_force[ 946] <= 8'h68;
  filter_in_data_log_force[ 947] <= 8'h68;
  filter_in_data_log_force[ 948] <= 8'h68;
  filter_in_data_log_force[ 949] <= 8'h68;
  filter_in_data_log_force[ 950] <= 8'h69;
  filter_in_data_log_force[ 951] <= 8'h69;
  filter_in_data_log_force[ 952] <= 8'h69;
  filter_in_data_log_force[ 953] <= 8'h69;
  filter_in_data_log_force[ 954] <= 8'h6a;
  filter_in_data_log_force[ 955] <= 8'h6a;
  filter_in_data_log_force[ 956] <= 8'h6a;
  filter_in_data_log_force[ 957] <= 8'h6a;
  filter_in_data_log_force[ 958] <= 8'h6b;
  filter_in_data_log_force[ 959] <= 8'h6b;
  filter_in_data_log_force[ 960] <= 8'h6b;
  filter_in_data_log_force[ 961] <= 8'h6b;
  filter_in_data_log_force[ 962] <= 8'h6c;
  filter_in_data_log_force[ 963] <= 8'h6c;
  filter_in_data_log_force[ 964] <= 8'h6c;
  filter_in_data_log_force[ 965] <= 8'h6c;
  filter_in_data_log_force[ 966] <= 8'h6d;
  filter_in_data_log_force[ 967] <= 8'h6d;
  filter_in_data_log_force[ 968] <= 8'h6d;
  filter_in_data_log_force[ 969] <= 8'h6d;
  filter_in_data_log_force[ 970] <= 8'h6e;
  filter_in_data_log_force[ 971] <= 8'h6e;
  filter_in_data_log_force[ 972] <= 8'h6e;
  filter_in_data_log_force[ 973] <= 8'h6e;
  filter_in_data_log_force[ 974] <= 8'h6f;
  filter_in_data_log_force[ 975] <= 8'h6f;
  filter_in_data_log_force[ 976] <= 8'h6f;
  filter_in_data_log_force[ 977] <= 8'h6f;
  filter_in_data_log_force[ 978] <= 8'h70;
  filter_in_data_log_force[ 979] <= 8'h70;
  filter_in_data_log_force[ 980] <= 8'h70;
  filter_in_data_log_force[ 981] <= 8'h70;
  filter_in_data_log_force[ 982] <= 8'h71;
  filter_in_data_log_force[ 983] <= 8'h71;
  filter_in_data_log_force[ 984] <= 8'h71;
  filter_in_data_log_force[ 985] <= 8'h71;
  filter_in_data_log_force[ 986] <= 8'h72;
  filter_in_data_log_force[ 987] <= 8'h72;
  filter_in_data_log_force[ 988] <= 8'h72;
  filter_in_data_log_force[ 989] <= 8'h72;
  filter_in_data_log_force[ 990] <= 8'h73;
  filter_in_data_log_force[ 991] <= 8'h73;
  filter_in_data_log_force[ 992] <= 8'h73;
  filter_in_data_log_force[ 993] <= 8'h73;
  filter_in_data_log_force[ 994] <= 8'h74;
  filter_in_data_log_force[ 995] <= 8'h74;
  filter_in_data_log_force[ 996] <= 8'h74;
  filter_in_data_log_force[ 997] <= 8'h74;
  filter_in_data_log_force[ 998] <= 8'h75;
  filter_in_data_log_force[ 999] <= 8'h75;
  filter_in_data_log_force[1000] <= 8'h75;
  filter_in_data_log_force[1001] <= 8'h75;
  filter_in_data_log_force[1002] <= 8'h76;
  filter_in_data_log_force[1003] <= 8'h76;
  filter_in_data_log_force[1004] <= 8'h76;
  filter_in_data_log_force[1005] <= 8'h76;
  filter_in_data_log_force[1006] <= 8'h77;
  filter_in_data_log_force[1007] <= 8'h77;
  filter_in_data_log_force[1008] <= 8'h77;
  filter_in_data_log_force[1009] <= 8'h77;
  filter_in_data_log_force[1010] <= 8'h78;
  filter_in_data_log_force[1011] <= 8'h78;
  filter_in_data_log_force[1012] <= 8'h78;
  filter_in_data_log_force[1013] <= 8'h78;
  filter_in_data_log_force[1014] <= 8'h79;
  filter_in_data_log_force[1015] <= 8'h79;
  filter_in_data_log_force[1016] <= 8'h79;
  filter_in_data_log_force[1017] <= 8'h79;
  filter_in_data_log_force[1018] <= 8'h7a;
  filter_in_data_log_force[1019] <= 8'h7a;
  filter_in_data_log_force[1020] <= 8'h7a;
  filter_in_data_log_force[1021] <= 8'h7a;
  filter_in_data_log_force[1022] <= 8'h7b;
  filter_in_data_log_force[1023] <= 8'h7b;
  filter_in_data_log_force[1024] <= 8'h7b;
  filter_in_data_log_force[1025] <= 8'h7b;
  filter_in_data_log_force[1026] <= 8'h7c;
  filter_in_data_log_force[1027] <= 8'h7c;
  filter_in_data_log_force[1028] <= 8'h7c;
  filter_in_data_log_force[1029] <= 8'h7c;
  filter_in_data_log_force[1030] <= 8'h7d;
  filter_in_data_log_force[1031] <= 8'h7d;
  filter_in_data_log_force[1032] <= 8'h7d;
  filter_in_data_log_force[1033] <= 8'h7d;
  filter_in_data_log_force[1034] <= 8'h7e;
  filter_in_data_log_force[1035] <= 8'h7e;
  filter_in_data_log_force[1036] <= 8'h7e;
  filter_in_data_log_force[1037] <= 8'h7e;
  filter_in_data_log_force[1038] <= 8'h7f;
  filter_in_data_log_force[1039] <= 8'h7f;
  filter_in_data_log_force[1040] <= 8'h7f;
  filter_in_data_log_force[1041] <= 8'h7f;
  filter_in_data_log_force[1042] <= 8'h7f;
  filter_in_data_log_force[1043] <= 8'h7f;
  filter_in_data_log_force[1044] <= 8'h00;
  filter_in_data_log_force[1045] <= 8'h00;
  filter_in_data_log_force[1046] <= 8'h00;
  filter_in_data_log_force[1047] <= 8'h00;
  filter_in_data_log_force[1048] <= 8'h00;
  filter_in_data_log_force[1049] <= 8'h7f;
  filter_in_data_log_force[1050] <= 8'h7f;
  filter_in_data_log_force[1051] <= 8'h7f;
  filter_in_data_log_force[1052] <= 8'h7f;
  filter_in_data_log_force[1053] <= 8'h7f;
  filter_in_data_log_force[1054] <= 8'h7f;
  filter_in_data_log_force[1055] <= 8'h7f;
  filter_in_data_log_force[1056] <= 8'h7f;
  filter_in_data_log_force[1057] <= 8'h7f;
  filter_in_data_log_force[1058] <= 8'h7f;
  filter_in_data_log_force[1059] <= 8'h7f;
  filter_in_data_log_force[1060] <= 8'h7e;
  filter_in_data_log_force[1061] <= 8'h7d;
  filter_in_data_log_force[1062] <= 8'h7c;
  filter_in_data_log_force[1063] <= 8'h7a;
  filter_in_data_log_force[1064] <= 8'h79;
  filter_in_data_log_force[1065] <= 8'h77;
  filter_in_data_log_force[1066] <= 8'h74;
  filter_in_data_log_force[1067] <= 8'h71;
  filter_in_data_log_force[1068] <= 8'h6e;
  filter_in_data_log_force[1069] <= 8'h6a;
  filter_in_data_log_force[1070] <= 8'h65;
  filter_in_data_log_force[1071] <= 8'h60;
  filter_in_data_log_force[1072] <= 8'h5a;
  filter_in_data_log_force[1073] <= 8'h53;
  filter_in_data_log_force[1074] <= 8'h4b;
  filter_in_data_log_force[1075] <= 8'h43;
  filter_in_data_log_force[1076] <= 8'h3a;
  filter_in_data_log_force[1077] <= 8'h31;
  filter_in_data_log_force[1078] <= 8'h26;
  filter_in_data_log_force[1079] <= 8'h1b;
  filter_in_data_log_force[1080] <= 8'h10;
  filter_in_data_log_force[1081] <= 8'h04;
  filter_in_data_log_force[1082] <= 8'hf7;
  filter_in_data_log_force[1083] <= 8'heb;
  filter_in_data_log_force[1084] <= 8'hde;
  filter_in_data_log_force[1085] <= 8'hd1;
  filter_in_data_log_force[1086] <= 8'hc4;
  filter_in_data_log_force[1087] <= 8'hb8;
  filter_in_data_log_force[1088] <= 8'hac;
  filter_in_data_log_force[1089] <= 8'ha1;
  filter_in_data_log_force[1090] <= 8'h97;
  filter_in_data_log_force[1091] <= 8'h8f;
  filter_in_data_log_force[1092] <= 8'h88;
  filter_in_data_log_force[1093] <= 8'h83;
  filter_in_data_log_force[1094] <= 8'h81;
  filter_in_data_log_force[1095] <= 8'h80;
  filter_in_data_log_force[1096] <= 8'h82;
  filter_in_data_log_force[1097] <= 8'h87;
  filter_in_data_log_force[1098] <= 8'h8e;
  filter_in_data_log_force[1099] <= 8'h98;
  filter_in_data_log_force[1100] <= 8'ha4;
  filter_in_data_log_force[1101] <= 8'hb3;
  filter_in_data_log_force[1102] <= 8'hc4;
  filter_in_data_log_force[1103] <= 8'hd7;
  filter_in_data_log_force[1104] <= 8'hec;
  filter_in_data_log_force[1105] <= 8'h01;
  filter_in_data_log_force[1106] <= 8'h16;
  filter_in_data_log_force[1107] <= 8'h2c;
  filter_in_data_log_force[1108] <= 8'h40;
  filter_in_data_log_force[1109] <= 8'h53;
  filter_in_data_log_force[1110] <= 8'h63;
  filter_in_data_log_force[1111] <= 8'h70;
  filter_in_data_log_force[1112] <= 8'h7a;
  filter_in_data_log_force[1113] <= 8'h7f;
  filter_in_data_log_force[1114] <= 8'h7f;
  filter_in_data_log_force[1115] <= 8'h7b;
  filter_in_data_log_force[1116] <= 8'h72;
  filter_in_data_log_force[1117] <= 8'h64;
  filter_in_data_log_force[1118] <= 8'h51;
  filter_in_data_log_force[1119] <= 8'h3b;
  filter_in_data_log_force[1120] <= 8'h22;
  filter_in_data_log_force[1121] <= 8'h07;
  filter_in_data_log_force[1122] <= 8'heb;
  filter_in_data_log_force[1123] <= 8'hd0;
  filter_in_data_log_force[1124] <= 8'hb7;
  filter_in_data_log_force[1125] <= 8'ha1;
  filter_in_data_log_force[1126] <= 8'h90;
  filter_in_data_log_force[1127] <= 8'h85;
  filter_in_data_log_force[1128] <= 8'h80;
  filter_in_data_log_force[1129] <= 8'h83;
  filter_in_data_log_force[1130] <= 8'h8d;
  filter_in_data_log_force[1131] <= 8'h9e;
  filter_in_data_log_force[1132] <= 8'hb5;
  filter_in_data_log_force[1133] <= 8'hd1;
  filter_in_data_log_force[1134] <= 8'hf0;
  filter_in_data_log_force[1135] <= 8'h11;
  filter_in_data_log_force[1136] <= 8'h31;
  filter_in_data_log_force[1137] <= 8'h4e;
  filter_in_data_log_force[1138] <= 8'h66;
  filter_in_data_log_force[1139] <= 8'h77;
  filter_in_data_log_force[1140] <= 8'h7f;
  filter_in_data_log_force[1141] <= 8'h7e;
  filter_in_data_log_force[1142] <= 8'h73;
  filter_in_data_log_force[1143] <= 8'h5f;
  filter_in_data_log_force[1144] <= 8'h44;
  filter_in_data_log_force[1145] <= 8'h22;
  filter_in_data_log_force[1146] <= 8'hfd;
  filter_in_data_log_force[1147] <= 8'hd8;
  filter_in_data_log_force[1148] <= 8'hb7;
  filter_in_data_log_force[1149] <= 8'h9b;
  filter_in_data_log_force[1150] <= 8'h88;
  filter_in_data_log_force[1151] <= 8'h80;
  filter_in_data_log_force[1152] <= 8'h84;
  filter_in_data_log_force[1153] <= 8'h94;
  filter_in_data_log_force[1154] <= 8'haf;
  filter_in_data_log_force[1155] <= 8'hd2;
  filter_in_data_log_force[1156] <= 8'hfa;
  filter_in_data_log_force[1157] <= 8'h22;
  filter_in_data_log_force[1158] <= 8'h48;
  filter_in_data_log_force[1159] <= 8'h67;
  filter_in_data_log_force[1160] <= 8'h7a;
  filter_in_data_log_force[1161] <= 8'h7f;
  filter_in_data_log_force[1162] <= 8'h78;
  filter_in_data_log_force[1163] <= 8'h61;
  filter_in_data_log_force[1164] <= 8'h40;
  filter_in_data_log_force[1165] <= 8'h16;
  filter_in_data_log_force[1166] <= 8'he9;
  filter_in_data_log_force[1167] <= 8'hbf;
  filter_in_data_log_force[1168] <= 8'h9d;
  filter_in_data_log_force[1169] <= 8'h87;
  filter_in_data_log_force[1170] <= 8'h80;
  filter_in_data_log_force[1171] <= 8'h8a;
  filter_in_data_log_force[1172] <= 8'ha5;
  filter_in_data_log_force[1173] <= 8'hcb;
  filter_in_data_log_force[1174] <= 8'hfa;
  filter_in_data_log_force[1175] <= 8'h29;
  filter_in_data_log_force[1176] <= 8'h53;
  filter_in_data_log_force[1177] <= 8'h72;
  filter_in_data_log_force[1178] <= 8'h7f;
  filter_in_data_log_force[1179] <= 8'h7a;
  filter_in_data_log_force[1180] <= 8'h63;
  filter_in_data_log_force[1181] <= 8'h3c;
  filter_in_data_log_force[1182] <= 8'h0b;
  filter_in_data_log_force[1183] <= 8'hd8;
  filter_in_data_log_force[1184] <= 8'hac;
  filter_in_data_log_force[1185] <= 8'h8c;
  filter_in_data_log_force[1186] <= 8'h80;
  filter_in_data_log_force[1187] <= 8'h89;
  filter_in_data_log_force[1188] <= 8'ha7;
  filter_in_data_log_force[1189] <= 8'hd4;
  filter_in_data_log_force[1190] <= 8'h09;
  filter_in_data_log_force[1191] <= 8'h3d;
  filter_in_data_log_force[1192] <= 8'h66;
  filter_in_data_log_force[1193] <= 8'h7d;
  filter_in_data_log_force[1194] <= 8'h7d;
  filter_in_data_log_force[1195] <= 8'h65;
  filter_in_data_log_force[1196] <= 8'h3a;
  filter_in_data_log_force[1197] <= 8'h03;
  filter_in_data_log_force[1198] <= 8'hcc;
  filter_in_data_log_force[1199] <= 8'h9e;
  filter_in_data_log_force[1200] <= 8'h84;
  filter_in_data_log_force[1201] <= 8'h83;
  filter_in_data_log_force[1202] <= 8'h9b;
  filter_in_data_log_force[1203] <= 8'hc9;
  filter_in_data_log_force[1204] <= 8'h03;
  filter_in_data_log_force[1205] <= 8'h3c;
  filter_in_data_log_force[1206] <= 8'h69;
  filter_in_data_log_force[1207] <= 8'h7f;
  filter_in_data_log_force[1208] <= 8'h79;
  filter_in_data_log_force[1209] <= 8'h57;
  filter_in_data_log_force[1210] <= 8'h21;
  filter_in_data_log_force[1211] <= 8'he4;
  filter_in_data_log_force[1212] <= 8'had;
  filter_in_data_log_force[1213] <= 8'h89;
  filter_in_data_log_force[1214] <= 8'h81;
  filter_in_data_log_force[1215] <= 8'h98;
  filter_in_data_log_force[1216] <= 8'hc9;
  filter_in_data_log_force[1217] <= 8'h08;
  filter_in_data_log_force[1218] <= 8'h45;
  filter_in_data_log_force[1219] <= 8'h71;
  filter_in_data_log_force[1220] <= 8'h7f;
  filter_in_data_log_force[1221] <= 8'h6e;
  filter_in_data_log_force[1222] <= 8'h3f;
  filter_in_data_log_force[1223] <= 8'hff;
  filter_in_data_log_force[1224] <= 8'hbf;
  filter_in_data_log_force[1225] <= 8'h90;
  filter_in_data_log_force[1226] <= 8'h80;
  filter_in_data_log_force[1227] <= 8'h93;
  filter_in_data_log_force[1228] <= 8'hc5;
  filter_in_data_log_force[1229] <= 8'h08;
  filter_in_data_log_force[1230] <= 8'h49;
  filter_in_data_log_force[1231] <= 8'h75;
  filter_in_data_log_force[1232] <= 8'h7f;
  filter_in_data_log_force[1233] <= 8'h64;
  filter_in_data_log_force[1234] <= 8'h2a;
  filter_in_data_log_force[1235] <= 8'he4;
  filter_in_data_log_force[1236] <= 8'ha6;
  filter_in_data_log_force[1237] <= 8'h83;
  filter_in_data_log_force[1238] <= 8'h88;
  filter_in_data_log_force[1239] <= 8'hb2;
  filter_in_data_log_force[1240] <= 8'hf5;
  filter_in_data_log_force[1241] <= 8'h3d;
  filter_in_data_log_force[1242] <= 8'h70;
  filter_in_data_log_force[1243] <= 8'h7f;
  filter_in_data_log_force[1244] <= 8'h64;
  filter_in_data_log_force[1245] <= 8'h27;
  filter_in_data_log_force[1246] <= 8'hdd;
  filter_in_data_log_force[1247] <= 8'h9e;
  filter_in_data_log_force[1248] <= 8'h81;
  filter_in_data_log_force[1249] <= 8'h90;
  filter_in_data_log_force[1250] <= 8'hc6;
  filter_in_data_log_force[1251] <= 8'h12;
  filter_in_data_log_force[1252] <= 8'h57;
  filter_in_data_log_force[1253] <= 8'h7d;
  filter_in_data_log_force[1254] <= 8'h76;
  filter_in_data_log_force[1255] <= 8'h42;
  filter_in_data_log_force[1256] <= 8'hf6;
  filter_in_data_log_force[1257] <= 8'hae;
  filter_in_data_log_force[1258] <= 8'h84;
  filter_in_data_log_force[1259] <= 8'h89;
  filter_in_data_log_force[1260] <= 8'hbd;
  filter_in_data_log_force[1261] <= 8'h0b;
  filter_in_data_log_force[1262] <= 8'h55;
  filter_in_data_log_force[1263] <= 8'h7d;
  filter_in_data_log_force[1264] <= 8'h74;
  filter_in_data_log_force[1265] <= 8'h3b;
  filter_in_data_log_force[1266] <= 8'hea;
  filter_in_data_log_force[1267] <= 8'ha2;
  filter_in_data_log_force[1268] <= 8'h80;
  filter_in_data_log_force[1269] <= 8'h95;
  filter_in_data_log_force[1270] <= 8'hd6;
  filter_in_data_log_force[1271] <= 8'h2a;
  filter_in_data_log_force[1272] <= 8'h6c;
  filter_in_data_log_force[1273] <= 8'h7f;
  filter_in_data_log_force[1274] <= 8'h5b;
  filter_in_data_log_force[1275] <= 8'h0e;
  filter_in_data_log_force[1276] <= 8'hbb;
  filter_in_data_log_force[1277] <= 8'h86;
  filter_in_data_log_force[1278] <= 8'h89;
  filter_in_data_log_force[1279] <= 8'hc2;
  filter_in_data_log_force[1280] <= 8'h18;
  filter_in_data_log_force[1281] <= 8'h63;
  filter_in_data_log_force[1282] <= 8'h7f;
  filter_in_data_log_force[1283] <= 8'h61;
  filter_in_data_log_force[1284] <= 8'h13;
  filter_in_data_log_force[1285] <= 8'hbc;
  filter_in_data_log_force[1286] <= 8'h86;
  filter_in_data_log_force[1287] <= 8'h8b;
  filter_in_data_log_force[1288] <= 8'hca;
  filter_in_data_log_force[1289] <= 8'h23;
  filter_in_data_log_force[1290] <= 8'h6c;
  filter_in_data_log_force[1291] <= 8'h7e;
  filter_in_data_log_force[1292] <= 8'h51;
  filter_in_data_log_force[1293] <= 8'hf9;
  filter_in_data_log_force[1294] <= 8'ha5;
  filter_in_data_log_force[1295] <= 8'h80;
  filter_in_data_log_force[1296] <= 8'h9e;
  filter_in_data_log_force[1297] <= 8'hf0;
  filter_in_data_log_force[1298] <= 8'h4a;
  filter_in_data_log_force[1299] <= 8'h7d;
  filter_in_data_log_force[1300] <= 8'h6d;
  filter_in_data_log_force[1301] <= 8'h21;
  filter_in_data_log_force[1302] <= 8'hc3;
  filter_in_data_log_force[1303] <= 8'h86;
  filter_in_data_log_force[1304] <= 8'h8d;
  filter_in_data_log_force[1305] <= 8'hd5;
  filter_in_data_log_force[1306] <= 8'h35;
  filter_in_data_log_force[1307] <= 8'h77;
  filter_in_data_log_force[1308] <= 8'h75;
  filter_in_data_log_force[1309] <= 8'h2f;
  filter_in_data_log_force[1310] <= 8'hce;
  filter_in_data_log_force[1311] <= 8'h89;
  filter_in_data_log_force[1312] <= 8'h8b;
  filter_in_data_log_force[1313] <= 8'hd2;
  filter_in_data_log_force[1314] <= 8'h35;
  filter_in_data_log_force[1315] <= 8'h79;
  filter_in_data_log_force[1316] <= 8'h73;
  filter_in_data_log_force[1317] <= 8'h27;
  filter_in_data_log_force[1318] <= 8'hc2;
  filter_in_data_log_force[1319] <= 8'h84;
  filter_in_data_log_force[1320] <= 8'h93;
  filter_in_data_log_force[1321] <= 8'he7;
  filter_in_data_log_force[1322] <= 8'h4b;
  filter_in_data_log_force[1323] <= 8'h7f;
  filter_in_data_log_force[1324] <= 8'h62;
  filter_in_data_log_force[1325] <= 8'h05;
  filter_in_data_log_force[1326] <= 8'ha5;
  filter_in_data_log_force[1327] <= 8'h80;
  filter_in_data_log_force[1328] <= 8'hb0;
  filter_in_data_log_force[1329] <= 8'h15;
  filter_in_data_log_force[1330] <= 8'h6c;
  filter_in_data_log_force[1331] <= 8'h7b;
  filter_in_data_log_force[1332] <= 8'h36;
  filter_in_data_log_force[1333] <= 8'hcc;
  filter_in_data_log_force[1334] <= 8'h86;
  filter_in_data_log_force[1335] <= 8'h94;
  filter_in_data_log_force[1336] <= 8'hed;
  filter_in_data_log_force[1337] <= 8'h54;
  filter_in_data_log_force[1338] <= 8'h7f;
  filter_in_data_log_force[1339] <= 8'h51;
  filter_in_data_log_force[1340] <= 8'he8;
  filter_in_data_log_force[1341] <= 8'h90;
  filter_in_data_log_force[1342] <= 8'h89;
  filter_in_data_log_force[1343] <= 8'hd9;
  filter_in_data_log_force[1344] <= 8'h46;
  filter_in_data_log_force[1345] <= 8'h7f;
  filter_in_data_log_force[1346] <= 8'h5a;
  filter_in_data_log_force[1347] <= 8'hf2;
  filter_in_data_log_force[1348] <= 8'h94;
  filter_in_data_log_force[1349] <= 8'h87;
  filter_in_data_log_force[1350] <= 8'hd7;
  filter_in_data_log_force[1351] <= 8'h46;
  filter_in_data_log_force[1352] <= 8'h7f;
  filter_in_data_log_force[1353] <= 8'h56;
  filter_in_data_log_force[1354] <= 8'he9;
  filter_in_data_log_force[1355] <= 8'h8e;
  filter_in_data_log_force[1356] <= 8'h8d;
  filter_in_data_log_force[1357] <= 8'he7;
  filter_in_data_log_force[1358] <= 8'h56;
  filter_in_data_log_force[1359] <= 8'h7f;
  filter_in_data_log_force[1360] <= 8'h42;
  filter_in_data_log_force[1361] <= 8'hcf;
  filter_in_data_log_force[1362] <= 8'h83;
  filter_in_data_log_force[1363] <= 8'h9f;
  filter_in_data_log_force[1364] <= 8'h0b;
  filter_in_data_log_force[1365] <= 8'h6e;
  filter_in_data_log_force[1366] <= 8'h75;
  filter_in_data_log_force[1367] <= 8'h19;
  filter_in_data_log_force[1368] <= 8'ha8;
  filter_in_data_log_force[1369] <= 8'h81;
  filter_in_data_log_force[1370] <= 8'hc8;
  filter_in_data_log_force[1371] <= 8'h3f;
  filter_in_data_log_force[1372] <= 8'h7f;
  filter_in_data_log_force[1373] <= 8'h51;
  filter_in_data_log_force[1374] <= 8'hdb;
  filter_in_data_log_force[1375] <= 8'h86;
  filter_in_data_log_force[1376] <= 8'h9d;
  filter_in_data_log_force[1377] <= 8'h0c;
  filter_in_data_log_force[1378] <= 8'h71;
  filter_in_data_log_force[1379] <= 8'h70;
  filter_in_data_log_force[1380] <= 8'h09;
  filter_in_data_log_force[1381] <= 8'h9a;
  filter_in_data_log_force[1382] <= 8'h88;
  filter_in_data_log_force[1383] <= 8'he5;
  filter_in_data_log_force[1384] <= 8'h5c;
  filter_in_data_log_force[1385] <= 8'h7c;
  filter_in_data_log_force[1386] <= 8'h28;
  filter_in_data_log_force[1387] <= 8'hae;
  filter_in_data_log_force[1388] <= 8'h81;
  filter_in_data_log_force[1389] <= 8'hcd;
  filter_in_data_log_force[1390] <= 8'h4a;
  filter_in_data_log_force[1391] <= 8'h7f;
  filter_in_data_log_force[1392] <= 8'h39;
  filter_in_data_log_force[1393] <= 8'hbb;
  filter_in_data_log_force[1394] <= 8'h80;
  filter_in_data_log_force[1395] <= 8'hc3;
  filter_in_data_log_force[1396] <= 8'h43;
  filter_in_data_log_force[1397] <= 8'h7f;
  filter_in_data_log_force[1398] <= 8'h3d;
  filter_in_data_log_force[1399] <= 8'hbd;
  filter_in_data_log_force[1400] <= 8'h80;
  filter_in_data_log_force[1401] <= 8'hc5;
  filter_in_data_log_force[1402] <= 8'h46;
  filter_in_data_log_force[1403] <= 8'h7f;
  filter_in_data_log_force[1404] <= 8'h35;
  filter_in_data_log_force[1405] <= 8'hb3;
  filter_in_data_log_force[1406] <= 8'h81;
  filter_in_data_log_force[1407] <= 8'hd4;
  filter_in_data_log_force[1408] <= 8'h55;
  filter_in_data_log_force[1409] <= 8'h7c;
  filter_in_data_log_force[1410] <= 8'h1f;
  filter_in_data_log_force[1411] <= 8'ha1;
  filter_in_data_log_force[1412] <= 8'h88;
  filter_in_data_log_force[1413] <= 8'hf1;
  filter_in_data_log_force[1414] <= 8'h6a;
  filter_in_data_log_force[1415] <= 8'h70;
  filter_in_data_log_force[1416] <= 8'hfa;
  filter_in_data_log_force[1417] <= 8'h8b;
  filter_in_data_log_force[1418] <= 8'h9d;
  filter_in_data_log_force[1419] <= 8'h1d;
  filter_in_data_log_force[1420] <= 8'h7d;
  filter_in_data_log_force[1421] <= 8'h50;
  filter_in_data_log_force[1422] <= 8'hc9;
  filter_in_data_log_force[1423] <= 8'h80;
  filter_in_data_log_force[1424] <= 8'hc8;
  filter_in_data_log_force[1425] <= 8'h51;
  filter_in_data_log_force[1426] <= 8'h7c;
  filter_in_data_log_force[1427] <= 8'h18;
  filter_in_data_log_force[1428] <= 8'h98;
  filter_in_data_log_force[1429] <= 8'h91;
  filter_in_data_log_force[1430] <= 8'h0c;
  filter_in_data_log_force[1431] <= 8'h79;
  filter_in_data_log_force[1432] <= 8'h57;
  filter_in_data_log_force[1433] <= 8'hce;
  filter_in_data_log_force[1434] <= 8'h80;
  filter_in_data_log_force[1435] <= 8'hcc;
  filter_in_data_log_force[1436] <= 8'h57;
  filter_in_data_log_force[1437] <= 8'h79;
  filter_in_data_log_force[1438] <= 8'h08;
  filter_in_data_log_force[1439] <= 8'h8d;
  filter_in_data_log_force[1440] <= 8'h9f;
  filter_in_data_log_force[1441] <= 8'h29;
  filter_in_data_log_force[1442] <= 8'h7f;
  filter_in_data_log_force[1443] <= 8'h38;
  filter_in_data_log_force[1444] <= 8'haa;
  filter_in_data_log_force[1445] <= 8'h88;
  filter_in_data_log_force[1446] <= 8'hfd;
  filter_in_data_log_force[1447] <= 8'h76;
  filter_in_data_log_force[1448] <= 8'h59;
  filter_in_data_log_force[1449] <= 8'hca;
  filter_in_data_log_force[1450] <= 8'h80;
  filter_in_data_log_force[1451] <= 8'hdb;
  filter_in_data_log_force[1452] <= 8'h65;
  filter_in_data_log_force[1453] <= 8'h6d;
  filter_in_data_log_force[1454] <= 8'he6;
  filter_in_data_log_force[1455] <= 8'h81;
  filter_in_data_log_force[1456] <= 8'hc3;
  filter_in_data_log_force[1457] <= 8'h56;
  filter_in_data_log_force[1458] <= 8'h76;
  filter_in_data_log_force[1459] <= 8'hf9;
  filter_in_data_log_force[1460] <= 8'h85;
  filter_in_data_log_force[1461] <= 8'hb6;
  filter_in_data_log_force[1462] <= 8'h4b;
  filter_in_data_log_force[1463] <= 8'h7a;
  filter_in_data_log_force[1464] <= 8'h03;
  filter_in_data_log_force[1465] <= 8'h87;
  filter_in_data_log_force[1466] <= 8'hb2;
  filter_in_data_log_force[1467] <= 8'h48;
  filter_in_data_log_force[1468] <= 8'h7b;
  filter_in_data_log_force[1469] <= 8'h03;
  filter_in_data_log_force[1470] <= 8'h87;
  filter_in_data_log_force[1471] <= 8'hb5;
  filter_in_data_log_force[1472] <= 8'h4d;
  filter_in_data_log_force[1473] <= 8'h78;
  filter_in_data_log_force[1474] <= 8'hf9;
  filter_in_data_log_force[1475] <= 8'h84;
  filter_in_data_log_force[1476] <= 8'hc0;
  filter_in_data_log_force[1477] <= 8'h58;
  filter_in_data_log_force[1478] <= 8'h72;
  filter_in_data_log_force[1479] <= 8'he6;
  filter_in_data_log_force[1480] <= 8'h80;
  filter_in_data_log_force[1481] <= 8'hd5;
  filter_in_data_log_force[1482] <= 8'h69;
  filter_in_data_log_force[1483] <= 8'h63;
  filter_in_data_log_force[1484] <= 8'hcb;
  filter_in_data_log_force[1485] <= 8'h82;
  filter_in_data_log_force[1486] <= 8'hf4;
  filter_in_data_log_force[1487] <= 8'h78;
  filter_in_data_log_force[1488] <= 8'h48;
  filter_in_data_log_force[1489] <= 8'hab;
  filter_in_data_log_force[1490] <= 8'h8f;
  filter_in_data_log_force[1491] <= 8'h1e;
  filter_in_data_log_force[1492] <= 8'h7f;
  filter_in_data_log_force[1493] <= 8'h1e;
  filter_in_data_log_force[1494] <= 8'h8e;
  filter_in_data_log_force[1495] <= 8'hae;
  filter_in_data_log_force[1496] <= 8'h4d;
  filter_in_data_log_force[1497] <= 8'h75;
  filter_in_data_log_force[1498] <= 8'he7;
  filter_in_data_log_force[1499] <= 8'h80;
  filter_in_data_log_force[1500] <= 8'he2;
  filter_in_data_log_force[1501] <= 8'h74;
  filter_in_data_log_force[1502] <= 8'h4e;
  filter_in_data_log_force[1503] <= 8'had;
  filter_in_data_log_force[1504] <= 8'h90;
  filter_in_data_log_force[1505] <= 8'h27;
  filter_in_data_log_force[1506] <= 8'h7f;
  filter_in_data_log_force[1507] <= 8'h0b;
  filter_in_data_log_force[1508] <= 8'h85;
  filter_in_data_log_force[1509] <= 8'hc7;
  filter_in_data_log_force[1510] <= 8'h66;
  filter_in_data_log_force[1511] <= 8'h5e;
  filter_in_data_log_force[1512] <= 8'hbc;
  filter_in_data_log_force[1513] <= 8'h89;
  filter_in_data_log_force[1514] <= 8'h1b;
  filter_in_data_log_force[1515] <= 8'h7f;
  filter_in_data_log_force[1516] <= 8'h10;
  filter_in_data_log_force[1517] <= 8'h85;
  filter_in_data_log_force[1518] <= 8'hc9;
  filter_in_data_log_force[1519] <= 8'h69;
  filter_in_data_log_force[1520] <= 8'h58;
  filter_in_data_log_force[1521] <= 8'hb2;
  filter_in_data_log_force[1522] <= 8'h90;
  filter_in_data_log_force[1523] <= 8'h2e;
  filter_in_data_log_force[1524] <= 8'h7d;
  filter_in_data_log_force[1525] <= 8'hf6;
  filter_in_data_log_force[1526] <= 8'h80;
  filter_in_data_log_force[1527] <= 8'he8;
  filter_in_data_log_force[1528] <= 8'h7a;
  filter_in_data_log_force[1529] <= 8'h37;
  filter_in_data_log_force[1530] <= 8'h94;
  filter_in_data_log_force[1531] <= 8'hae;
  filter_in_data_log_force[1532] <= 8'h58;
  filter_in_data_log_force[1533] <= 8'h66;
  filter_in_data_log_force[1534] <= 8'hbf;
  filter_in_data_log_force[1535] <= 8'h8b;
  filter_in_data_log_force[1536] <= 8'h28;
  filter_in_data_log_force[1537] <= 8'h7d;
  filter_in_data_log_force[1538] <= 8'hf2;
  filter_in_data_log_force[1539] <= 8'h80;
  filter_in_data_log_force[1540] <= 8'hf5;
  filter_in_data_log_force[1541] <= 8'h7e;
  filter_in_data_log_force[1542] <= 8'h21;
  filter_in_data_log_force[1543] <= 8'h88;
  filter_in_data_log_force[1544] <= 8'hcb;
  filter_in_data_log_force[1545] <= 8'h70;
  filter_in_data_log_force[1546] <= 8'h47;
  filter_in_data_log_force[1547] <= 8'h9b;
  filter_in_data_log_force[1548] <= 8'hab;
  filter_in_data_log_force[1549] <= 8'h59;
  filter_in_data_log_force[1550] <= 8'h61;
  filter_in_data_log_force[1551] <= 8'hb3;
  filter_in_data_log_force[1552] <= 8'h95;
  filter_in_data_log_force[1553] <= 8'h41;
  filter_in_data_log_force[1554] <= 8'h72;
  filter_in_data_log_force[1555] <= 8'hcb;
  filter_in_data_log_force[1556] <= 8'h89;
  filter_in_data_log_force[1557] <= 8'h2b;
  filter_in_data_log_force[1558] <= 8'h7a;
  filter_in_data_log_force[1559] <= 8'hdf;
  filter_in_data_log_force[1560] <= 8'h83;
  filter_in_data_log_force[1561] <= 8'h19;
  filter_in_data_log_force[1562] <= 8'h7e;
  filter_in_data_log_force[1563] <= 8'hee;
  filter_in_data_log_force[1564] <= 8'h81;
  filter_in_data_log_force[1565] <= 8'h0d;
  filter_in_data_log_force[1566] <= 8'h7f;
  filter_in_data_log_force[1567] <= 8'hf7;
  filter_in_data_log_force[1568] <= 8'h80;
  filter_in_data_log_force[1569] <= 8'h07;
  filter_in_data_log_force[1570] <= 8'h7f;
  filter_in_data_log_force[1571] <= 8'hfa;
  filter_in_data_log_force[1572] <= 8'h80;
  filter_in_data_log_force[1573] <= 8'h07;
  filter_in_data_log_force[1574] <= 8'h7f;
  filter_in_data_log_force[1575] <= 8'hf7;
  filter_in_data_log_force[1576] <= 8'h80;
  filter_in_data_log_force[1577] <= 8'h0d;
  filter_in_data_log_force[1578] <= 8'h7f;
  filter_in_data_log_force[1579] <= 8'hed;
  filter_in_data_log_force[1580] <= 8'h82;
  filter_in_data_log_force[1581] <= 8'h19;
  filter_in_data_log_force[1582] <= 8'h7d;
  filter_in_data_log_force[1583] <= 8'hde;
  filter_in_data_log_force[1584] <= 8'h86;
  filter_in_data_log_force[1585] <= 8'h2b;
  filter_in_data_log_force[1586] <= 8'h76;
  filter_in_data_log_force[1587] <= 8'hca;
  filter_in_data_log_force[1588] <= 8'h8f;
  filter_in_data_log_force[1589] <= 8'h42;
  filter_in_data_log_force[1590] <= 8'h6a;
  filter_in_data_log_force[1591] <= 8'hb2;
  filter_in_data_log_force[1592] <= 8'h9f;
  filter_in_data_log_force[1593] <= 8'h5a;
  filter_in_data_log_force[1594] <= 8'h55;
  filter_in_data_log_force[1595] <= 8'h9a;
  filter_in_data_log_force[1596] <= 8'hba;
  filter_in_data_log_force[1597] <= 8'h70;
  filter_in_data_log_force[1598] <= 8'h34;
  filter_in_data_log_force[1599] <= 8'h87;
  filter_in_data_log_force[1600] <= 8'he0;
  filter_in_data_log_force[1601] <= 8'h7e;
  filter_in_data_log_force[1602] <= 8'h09;
  filter_in_data_log_force[1603] <= 8'h80;
  filter_in_data_log_force[1604] <= 8'h10;
  filter_in_data_log_force[1605] <= 8'h7d;
  filter_in_data_log_force[1606] <= 8'hd7;
  filter_in_data_log_force[1607] <= 8'h8c;
  filter_in_data_log_force[1608] <= 8'h42;
  filter_in_data_log_force[1609] <= 8'h65;
  filter_in_data_log_force[1610] <= 8'ha7;
  filter_in_data_log_force[1611] <= 8'hb0;
  filter_in_data_log_force[1612] <= 8'h6d;
  filter_in_data_log_force[1613] <= 8'h36;
  filter_in_data_log_force[1614] <= 8'h86;
  filter_in_data_log_force[1615] <= 8'hea;
  filter_in_data_log_force[1616] <= 8'h7f;
  filter_in_data_log_force[1617] <= 8'hf3;
  filter_in_data_log_force[1618] <= 8'h84;
  filter_in_data_log_force[1619] <= 8'h30;
  filter_in_data_log_force[1620] <= 8'h6f;
  filter_in_data_log_force[1621] <= 8'hb0;
  filter_in_data_log_force[1622] <= 8'haa;
  filter_in_data_log_force[1623] <= 8'h6b;
  filter_in_data_log_force[1624] <= 8'h35;
  filter_in_data_log_force[1625] <= 8'h85;
  filter_in_data_log_force[1626] <= 8'hf3;
  filter_in_data_log_force[1627] <= 8'h7f;
  filter_in_data_log_force[1628] <= 8'he2;
  filter_in_data_log_force[1629] <= 8'h8b;
  filter_in_data_log_force[1630] <= 8'h47;
  filter_in_data_log_force[1631] <= 8'h5c;
  filter_in_data_log_force[1632] <= 8'h98;
  filter_in_data_log_force[1633] <= 8'hca;
  filter_in_data_log_force[1634] <= 8'h7c;
  filter_in_data_log_force[1635] <= 8'h08;
  filter_in_data_log_force[1636] <= 8'h81;
  filter_in_data_log_force[1637] <= 8'h2a;
  filter_in_data_log_force[1638] <= 8'h6e;
  filter_in_data_log_force[1639] <= 8'haa;
  filter_in_data_log_force[1640] <= 8'hb5;
  filter_in_data_log_force[1641] <= 8'h75;
  filter_in_data_log_force[1642] <= 8'h1a;
  filter_in_data_log_force[1643] <= 8'h80;
  filter_in_data_log_force[1644] <= 8'h1d;
  filter_in_data_log_force[1645] <= 8'h73;
  filter_in_data_log_force[1646] <= 8'hb0;
  filter_in_data_log_force[1647] <= 8'hb0;
  filter_in_data_log_force[1648] <= 8'h74;
  filter_in_data_log_force[1649] <= 8'h1a;
  filter_in_data_log_force[1650] <= 8'h80;
  filter_in_data_log_force[1651] <= 8'h22;
  filter_in_data_log_force[1652] <= 8'h70;
  filter_in_data_log_force[1653] <= 8'ha8;
  filter_in_data_log_force[1654] <= 8'hbb;
  filter_in_data_log_force[1655] <= 8'h7a;
  filter_in_data_log_force[1656] <= 8'h08;
  filter_in_data_log_force[1657] <= 8'h82;
  filter_in_data_log_force[1658] <= 8'h39;
  filter_in_data_log_force[1659] <= 8'h60;
  filter_in_data_log_force[1660] <= 8'h95;
  filter_in_data_log_force[1661] <= 8'hd9;
  filter_in_data_log_force[1662] <= 8'h7f;
  filter_in_data_log_force[1663] <= 8'he2;
  filter_in_data_log_force[1664] <= 8'h91;
  filter_in_data_log_force[1665] <= 8'h5b;
  filter_in_data_log_force[1666] <= 8'h3c;
  filter_in_data_log_force[1667] <= 8'h83;
  filter_in_data_log_force[1668] <= 8'h0b;
  filter_in_data_log_force[1669] <= 8'h77;
  filter_in_data_log_force[1670] <= 8'hb0;
  filter_in_data_log_force[1671] <= 8'hb8;
  filter_in_data_log_force[1672] <= 8'h7b;
  filter_in_data_log_force[1673] <= 8'hfe;
  filter_in_data_log_force[1674] <= 8'h87;
  filter_in_data_log_force[1675] <= 8'h4c;
  filter_in_data_log_force[1676] <= 8'h4b;
  filter_in_data_log_force[1677] <= 8'h86;
  filter_in_data_log_force[1678] <= 8'h02;
  filter_in_data_log_force[1679] <= 8'h79;
  filter_in_data_log_force[1680] <= 8'hb1;
  filter_in_data_log_force[1681] <= 8'hbb;
  filter_in_data_log_force[1682] <= 8'h7c;
  filter_in_data_log_force[1683] <= 8'hf4;
  filter_in_data_log_force[1684] <= 8'h8c;
  filter_in_data_log_force[1685] <= 8'h5a;
  filter_in_data_log_force[1686] <= 8'h38;
  filter_in_data_log_force[1687] <= 8'h81;
  filter_in_data_log_force[1688] <= 8'h1f;
  filter_in_data_log_force[1689] <= 8'h6a;
  filter_in_data_log_force[1690] <= 8'h97;
  filter_in_data_log_force[1691] <= 8'he0;
  filter_in_data_log_force[1692] <= 8'h7f;
  filter_in_data_log_force[1693] <= 8'hc5;
  filter_in_data_log_force[1694] <= 8'hab;
  filter_in_data_log_force[1695] <= 8'h78;
  filter_in_data_log_force[1696] <= 8'hfd;
  filter_in_data_log_force[1697] <= 8'h8a;
  filter_in_data_log_force[1698] <= 8'h5a;
  filter_in_data_log_force[1699] <= 8'h33;
  filter_in_data_log_force[1700] <= 8'h80;
  filter_in_data_log_force[1701] <= 8'h2e;
  filter_in_data_log_force[1702] <= 8'h5d;
  filter_in_data_log_force[1703] <= 8'h8b;
  filter_in_data_log_force[1704] <= 8'hfe;
  filter_in_data_log_force[1705] <= 8'h76;
  filter_in_data_log_force[1706] <= 8'ha5;
  filter_in_data_log_force[1707] <= 8'hd2;
  filter_in_data_log_force[1708] <= 8'h7f;
  filter_in_data_log_force[1709] <= 8'hc8;
  filter_in_data_log_force[1710] <= 8'hae;
  filter_in_data_log_force[1711] <= 8'h7b;
  filter_in_data_log_force[1712] <= 8'hed;
  filter_in_data_log_force[1713] <= 8'h94;
  filter_in_data_log_force[1714] <= 8'h6c;
  filter_in_data_log_force[1715] <= 8'h12;
  filter_in_data_log_force[1716] <= 8'h86;
  filter_in_data_log_force[1717] <= 8'h56;
  filter_in_data_log_force[1718] <= 8'h31;
  filter_in_data_log_force[1719] <= 8'h80;
  filter_in_data_log_force[1720] <= 8'h3d;
  filter_in_data_log_force[1721] <= 8'h4b;
  filter_in_data_log_force[1722] <= 8'h82;
  filter_in_data_log_force[1723] <= 8'h24;
  filter_in_data_log_force[1724] <= 8'h5e;
  filter_in_data_log_force[1725] <= 8'h88;
  filter_in_data_log_force[1726] <= 8'h0d;
  filter_in_data_log_force[1727] <= 8'h6c;
  filter_in_data_log_force[1728] <= 8'h92;
  filter_in_data_log_force[1729] <= 8'hf9;
  filter_in_data_log_force[1730] <= 8'h75;
  filter_in_data_log_force[1731] <= 8'h9c;
  filter_in_data_log_force[1732] <= 8'he8;
  filter_in_data_log_force[1733] <= 8'h7a;
  filter_in_data_log_force[1734] <= 8'ha5;
  filter_in_data_log_force[1735] <= 8'hdb;
  filter_in_data_log_force[1736] <= 8'h7d;
  filter_in_data_log_force[1737] <= 8'had;
  filter_in_data_log_force[1738] <= 8'hd2;
  filter_in_data_log_force[1739] <= 8'h7f;
  filter_in_data_log_force[1740] <= 8'hb3;
  filter_in_data_log_force[1741] <= 8'hcc;
  filter_in_data_log_force[1742] <= 8'h7f;
  filter_in_data_log_force[1743] <= 8'hb6;
  filter_in_data_log_force[1744] <= 8'hca;
  filter_in_data_log_force[1745] <= 8'h7f;
  filter_in_data_log_force[1746] <= 8'hb7;
  filter_in_data_log_force[1747] <= 8'hca;
  filter_in_data_log_force[1748] <= 8'h7f;
  filter_in_data_log_force[1749] <= 8'hb4;
  filter_in_data_log_force[1750] <= 8'hce;
  filter_in_data_log_force[1751] <= 8'h7f;
  filter_in_data_log_force[1752] <= 8'haf;
  filter_in_data_log_force[1753] <= 8'hd5;
  filter_in_data_log_force[1754] <= 8'h7d;
  filter_in_data_log_force[1755] <= 8'ha8;
  filter_in_data_log_force[1756] <= 8'he0;
  filter_in_data_log_force[1757] <= 8'h7a;
  filter_in_data_log_force[1758] <= 8'h9e;
  filter_in_data_log_force[1759] <= 8'hee;
  filter_in_data_log_force[1760] <= 8'h74;
  filter_in_data_log_force[1761] <= 8'h94;
  filter_in_data_log_force[1762] <= 8'h00;
  filter_in_data_log_force[1763] <= 8'h6b;
  filter_in_data_log_force[1764] <= 8'h8b;
  filter_in_data_log_force[1765] <= 8'h15;
  filter_in_data_log_force[1766] <= 8'h5d;
  filter_in_data_log_force[1767] <= 8'h83;
  filter_in_data_log_force[1768] <= 8'h2e;
  filter_in_data_log_force[1769] <= 8'h4a;
  filter_in_data_log_force[1770] <= 8'h80;
  filter_in_data_log_force[1771] <= 8'h47;
  filter_in_data_log_force[1772] <= 8'h30;
  filter_in_data_log_force[1773] <= 8'h83;
  filter_in_data_log_force[1774] <= 8'h5f;
  filter_in_data_log_force[1775] <= 8'h10;
  filter_in_data_log_force[1776] <= 8'h8f;
  filter_in_data_log_force[1777] <= 8'h73;
  filter_in_data_log_force[1778] <= 8'heb;
  filter_in_data_log_force[1779] <= 8'ha6;
  filter_in_data_log_force[1780] <= 8'h7e;
  filter_in_data_log_force[1781] <= 8'hc6;
  filter_in_data_log_force[1782] <= 8'hc7;
  filter_in_data_log_force[1783] <= 8'h7e;
  filter_in_data_log_force[1784] <= 8'ha3;
  filter_in_data_log_force[1785] <= 8'hf1;
  filter_in_data_log_force[1786] <= 8'h6e;
  filter_in_data_log_force[1787] <= 8'h8a;
  filter_in_data_log_force[1788] <= 8'h21;
  filter_in_data_log_force[1789] <= 8'h4e;
  filter_in_data_log_force[1790] <= 8'h80;
  filter_in_data_log_force[1791] <= 8'h4f;
  filter_in_data_log_force[1792] <= 8'h1f;
  filter_in_data_log_force[1793] <= 8'h8b;
  filter_in_data_log_force[1794] <= 8'h72;
  filter_in_data_log_force[1795] <= 8'he7;
  filter_in_data_log_force[1796] <= 8'had;
  filter_in_data_log_force[1797] <= 8'h7f;
  filter_in_data_log_force[1798] <= 8'hb1;
  filter_in_data_log_force[1799] <= 8'he3;
  filter_in_data_log_force[1800] <= 8'h73;
  filter_in_data_log_force[1801] <= 8'h8b;
  filter_in_data_log_force[1802] <= 8'h23;
  filter_in_data_log_force[1803] <= 8'h48;
  filter_in_data_log_force[1804] <= 8'h81;
  filter_in_data_log_force[1805] <= 8'h5c;
  filter_in_data_log_force[1806] <= 8'h08;
  filter_in_data_log_force[1807] <= 8'h9a;
  filter_in_data_log_force[1808] <= 8'h7d;
  filter_in_data_log_force[1809] <= 8'hc2;
  filter_in_data_log_force[1810] <= 8'hd4;
  filter_in_data_log_force[1811] <= 8'h77;
  filter_in_data_log_force[1812] <= 8'h8e;
  filter_in_data_log_force[1813] <= 8'h20;
  filter_in_data_log_force[1814] <= 8'h47;
  filter_in_data_log_force[1815] <= 8'h81;
  filter_in_data_log_force[1816] <= 8'h63;
  filter_in_data_log_force[1817] <= 8'hfa;
  filter_in_data_log_force[1818] <= 8'ha6;
  filter_in_data_log_force[1819] <= 8'h7f;
  filter_in_data_log_force[1820] <= 8'hac;
  filter_in_data_log_force[1821] <= 8'hf3;
  filter_in_data_log_force[1822] <= 8'h66;
  filter_in_data_log_force[1823] <= 8'h82;
  filter_in_data_log_force[1824] <= 8'h48;
  filter_in_data_log_force[1825] <= 8'h1b;
  filter_in_data_log_force[1826] <= 8'h93;
  filter_in_data_log_force[1827] <= 8'h7c;
  filter_in_data_log_force[1828] <= 8'hc0;
  filter_in_data_log_force[1829] <= 8'hde;
  filter_in_data_log_force[1830] <= 8'h70;
  filter_in_data_log_force[1831] <= 8'h85;
  filter_in_data_log_force[1832] <= 8'h3d;
  filter_in_data_log_force[1833] <= 8'h24;
  filter_in_data_log_force[1834] <= 8'h90;
  filter_in_data_log_force[1835] <= 8'h7b;
  filter_in_data_log_force[1836] <= 8'hc0;
  filter_in_data_log_force[1837] <= 8'he1;
  filter_in_data_log_force[1838] <= 8'h6d;
  filter_in_data_log_force[1839] <= 8'h83;
  filter_in_data_log_force[1840] <= 8'h48;
  filter_in_data_log_force[1841] <= 8'h14;
  filter_in_data_log_force[1842] <= 8'h9a;
  filter_in_data_log_force[1843] <= 8'h7f;
  filter_in_data_log_force[1844] <= 8'hac;
  filter_in_data_log_force[1845] <= 8'hfd;
  filter_in_data_log_force[1846] <= 8'h59;
  filter_in_data_log_force[1847] <= 8'h80;
  filter_in_data_log_force[1848] <= 8'h64;
  filter_in_data_log_force[1849] <= 8'hec;
  filter_in_data_log_force[1850] <= 8'hba;
  filter_in_data_log_force[1851] <= 8'h7c;
  filter_in_data_log_force[1852] <= 8'h8d;
  filter_in_data_log_force[1853] <= 8'h30;
  filter_in_data_log_force[1854] <= 8'h2a;
  filter_in_data_log_force[1855] <= 8'h91;
  filter_in_data_log_force[1856] <= 8'h7e;
  filter_in_data_log_force[1857] <= 8'hb1;
  filter_in_data_log_force[1858] <= 8'hfa;
  filter_in_data_log_force[1859] <= 8'h57;
  filter_in_data_log_force[1860] <= 8'h81;
  filter_in_data_log_force[1861] <= 8'h6b;
  filter_in_data_log_force[1862] <= 8'hdb;
  filter_in_data_log_force[1863] <= 8'hce;
  filter_in_data_log_force[1864] <= 8'h72;
  filter_in_data_log_force[1865] <= 8'h83;
  filter_in_data_log_force[1866] <= 8'h50;
  filter_in_data_log_force[1867] <= 8'h00;
  filter_in_data_log_force[1868] <= 8'haf;
  filter_in_data_log_force[1869] <= 8'h7d;
  filter_in_data_log_force[1870] <= 8'h8d;
  filter_in_data_log_force[1871] <= 8'h37;
  filter_in_data_log_force[1872] <= 8'h1c;
  filter_in_data_log_force[1873] <= 8'h9d;
  filter_in_data_log_force[1874] <= 8'h7f;
  filter_in_data_log_force[1875] <= 8'h99;
  filter_in_data_log_force[1876] <= 8'h24;
  filter_in_data_log_force[1877] <= 8'h2e;
  filter_in_data_log_force[1878] <= 8'h93;
  filter_in_data_log_force[1879] <= 8'h7f;
  filter_in_data_log_force[1880] <= 8'ha1;
  filter_in_data_log_force[1881] <= 8'h19;
  filter_in_data_log_force[1882] <= 8'h36;
  filter_in_data_log_force[1883] <= 8'h90;
  filter_in_data_log_force[1884] <= 8'h7f;
  filter_in_data_log_force[1885] <= 8'ha3;
  filter_in_data_log_force[1886] <= 8'h18;
  filter_in_data_log_force[1887] <= 8'h35;
  filter_in_data_log_force[1888] <= 8'h91;
  filter_in_data_log_force[1889] <= 8'h7f;
  filter_in_data_log_force[1890] <= 8'h9e;
  filter_in_data_log_force[1891] <= 8'h21;
  filter_in_data_log_force[1892] <= 8'h2c;
  filter_in_data_log_force[1893] <= 8'h98;
  filter_in_data_log_force[1894] <= 8'h7f;
  filter_in_data_log_force[1895] <= 8'h95;
  filter_in_data_log_force[1896] <= 8'h32;
  filter_in_data_log_force[1897] <= 8'h18;
  filter_in_data_log_force[1898] <= 8'ha6;
  filter_in_data_log_force[1899] <= 8'h7d;
  filter_in_data_log_force[1900] <= 8'h89;
  filter_in_data_log_force[1901] <= 8'h4a;
  filter_in_data_log_force[1902] <= 8'hfb;
  filter_in_data_log_force[1903] <= 8'hbf;
  filter_in_data_log_force[1904] <= 8'h72;
  filter_in_data_log_force[1905] <= 8'h81;
  filter_in_data_log_force[1906] <= 8'h65;
  filter_in_data_log_force[1907] <= 8'hd5;
  filter_in_data_log_force[1908] <= 8'he5;
  filter_in_data_log_force[1909] <= 8'h59;
  filter_in_data_log_force[1910] <= 8'h84;
  filter_in_data_log_force[1911] <= 8'h7a;
  filter_in_data_log_force[1912] <= 8'hab;
  filter_in_data_log_force[1913] <= 8'h18;
  filter_in_data_log_force[1914] <= 8'h2c;
  filter_in_data_log_force[1915] <= 8'h9c;
  filter_in_data_log_force[1916] <= 8'h7f;
  filter_in_data_log_force[1917] <= 8'h89;
  filter_in_data_log_force[1918] <= 8'h4e;
  filter_in_data_log_force[1919] <= 8'hef;
  filter_in_data_log_force[1920] <= 8'hd0;
  filter_in_data_log_force[1921] <= 8'h65;
  filter_in_data_log_force[1922] <= 8'h81;
  filter_in_data_log_force[1923] <= 8'h78;
  filter_in_data_log_force[1924] <= 8'hae;
  filter_in_data_log_force[1925] <= 8'h18;
  filter_in_data_log_force[1926] <= 8'h28;
  filter_in_data_log_force[1927] <= 8'ha3;
  filter_in_data_log_force[1928] <= 8'h7c;
  filter_in_data_log_force[1929] <= 8'h84;
  filter_in_data_log_force[1930] <= 8'h60;
  filter_in_data_log_force[1931] <= 8'hd4;
  filter_in_data_log_force[1932] <= 8'hef;
  filter_in_data_log_force[1933] <= 8'h4a;
  filter_in_data_log_force[1934] <= 8'h8e;
  filter_in_data_log_force[1935] <= 8'h7f;
  filter_in_data_log_force[1936] <= 8'h8e;
  filter_in_data_log_force[1937] <= 8'h4b;
  filter_in_data_log_force[1938] <= 8'hec;
  filter_in_data_log_force[1939] <= 8'hd9;
  filter_in_data_log_force[1940] <= 8'h59;
  filter_in_data_log_force[1941] <= 8'h88;
  filter_in_data_log_force[1942] <= 8'h7f;
  filter_in_data_log_force[1943] <= 8'h94;
  filter_in_data_log_force[1944] <= 8'h44;
  filter_in_data_log_force[1945] <= 8'hf2;
  filter_in_data_log_force[1946] <= 8'hd6;
  filter_in_data_log_force[1947] <= 8'h59;
  filter_in_data_log_force[1948] <= 8'h88;
  filter_in_data_log_force[1949] <= 8'h7f;
  filter_in_data_log_force[1950] <= 8'h90;
  filter_in_data_log_force[1951] <= 8'h4c;
  filter_in_data_log_force[1952] <= 8'he5;
  filter_in_data_log_force[1953] <= 8'he5;
  filter_in_data_log_force[1954] <= 8'h4b;
  filter_in_data_log_force[1955] <= 8'h91;
  filter_in_data_log_force[1956] <= 8'h7f;
  filter_in_data_log_force[1957] <= 8'h86;
  filter_in_data_log_force[1958] <= 8'h61;
  filter_in_data_log_force[1959] <= 8'hc7;
  filter_in_data_log_force[1960] <= 8'h07;
  filter_in_data_log_force[1961] <= 8'h2b;
  filter_in_data_log_force[1962] <= 8'haa;
  filter_in_data_log_force[1963] <= 8'h74;
  filter_in_data_log_force[1964] <= 8'h80;
  filter_in_data_log_force[1965] <= 8'h79;
  filter_in_data_log_force[1966] <= 8'h9f;
  filter_in_data_log_force[1967] <= 8'h3a;
  filter_in_data_log_force[1968] <= 8'hf4;
  filter_in_data_log_force[1969] <= 8'hdd;
  filter_in_data_log_force[1970] <= 8'h4d;
  filter_in_data_log_force[1971] <= 8'h93;
  filter_in_data_log_force[1972] <= 8'h7e;
  filter_in_data_log_force[1973] <= 8'h82;
  filter_in_data_log_force[1974] <= 8'h6e;
  filter_in_data_log_force[1975] <= 8'haf;
  filter_in_data_log_force[1976] <= 8'h29;
  filter_in_data_log_force[1977] <= 8'h03;
  filter_in_data_log_force[1978] <= 8'hd2;
  filter_in_data_log_force[1979] <= 8'h54;
  filter_in_data_log_force[1980] <= 8'h91;
  filter_in_data_log_force[1981] <= 8'h7e;
  filter_in_data_log_force[1982] <= 8'h82;
  filter_in_data_log_force[1983] <= 8'h71;
  filter_in_data_log_force[1984] <= 8'ha9;
  filter_in_data_log_force[1985] <= 8'h35;
  filter_in_data_log_force[1986] <= 8'hf3;
  filter_in_data_log_force[1987] <= 8'he4;
  filter_in_data_log_force[1988] <= 8'h41;
  filter_in_data_log_force[1989] <= 8'ha0;
  filter_in_data_log_force[1990] <= 8'h75;
  filter_in_data_log_force[1991] <= 8'h81;
  filter_in_data_log_force[1992] <= 8'h7d;
  filter_in_data_log_force[1993] <= 8'h90;
  filter_in_data_log_force[1994] <= 8'h59;
  filter_in_data_log_force[1995] <= 8'hc6;
  filter_in_data_log_force[1996] <= 8'h17;
  filter_in_data_log_force[1997] <= 8'h0e;
  filter_in_data_log_force[1998] <= 8'hce;
  filter_in_data_log_force[1999] <= 8'h51;
  filter_in_data_log_force[2000] <= 8'h97;
  filter_in_data_log_force[2001] <= 8'h79;
  filter_in_data_log_force[2002] <= 8'h80;
  filter_in_data_log_force[2003] <= 8'h7d;
  filter_in_data_log_force[2004] <= 8'h8f;
  filter_in_data_log_force[2005] <= 8'h5d;
  filter_in_data_log_force[2006] <= 8'hbd;
  filter_in_data_log_force[2007] <= 8'h25;
  filter_in_data_log_force[2008] <= 8'hfb;
  filter_in_data_log_force[2009] <= 8'he5;
  filter_in_data_log_force[2010] <= 8'h3a;
  filter_in_data_log_force[2011] <= 8'hac;
  filter_in_data_log_force[2012] <= 8'h69;
  filter_in_data_log_force[2013] <= 8'h89;
  filter_in_data_log_force[2014] <= 8'h7f;
  filter_in_data_log_force[2015] <= 8'h81;
  filter_in_data_log_force[2016] <= 8'h79;
  filter_in_data_log_force[2017] <= 8'h94;
  filter_in_data_log_force[2018] <= 8'h5a;
  filter_in_data_log_force[2019] <= 8'hbd;
  filter_in_data_log_force[2020] <= 8'h2a;
  filter_in_data_log_force[2021] <= 8'hf2;
  filter_in_data_log_force[2022] <= 8'hf3;
  filter_in_data_log_force[2023] <= 8'h28;
  filter_in_data_log_force[2024] <= 8'hc0;
  filter_in_data_log_force[2025] <= 8'h55;
  filter_in_data_log_force[2026] <= 8'h99;
  filter_in_data_log_force[2027] <= 8'h74;
  filter_in_data_log_force[2028] <= 8'h84;
  filter_in_data_log_force[2029] <= 8'h7f;
  filter_in_data_log_force[2030] <= 8'h81;
  filter_in_data_log_force[2031] <= 8'h79;
  filter_in_data_log_force[2032] <= 8'h91;
  filter_in_data_log_force[2033] <= 8'h62;
  filter_in_data_log_force[2034] <= 8'hae;
  filter_in_data_log_force[2035] <= 8'h40;
  filter_in_data_log_force[2036] <= 8'hd4;
  filter_in_data_log_force[2037] <= 8'h17;
  filter_in_data_log_force[2038] <= 8'hff;
  filter_in_data_log_force[2039] <= 8'hed;
  filter_in_data_log_force[2040] <= 8'h27;
  filter_in_data_log_force[2041] <= 8'hc6;
  filter_in_data_log_force[2042] <= 8'h4b;
  filter_in_data_log_force[2043] <= 8'ha6;
  filter_in_data_log_force[2044] <= 8'h66;
  filter_in_data_log_force[2045] <= 8'h90;
  filter_in_data_log_force[2046] <= 8'h78;
  filter_in_data_log_force[2047] <= 8'h83;
  filter_in_data_log_force[2048] <= 8'h7f;
  filter_in_data_log_force[2049] <= 8'h80;
  filter_in_data_log_force[2050] <= 8'h7e;
  filter_in_data_log_force[2051] <= 8'h86;
  filter_in_data_log_force[2052] <= 8'h74;
  filter_in_data_log_force[2053] <= 8'h93;
  filter_in_data_log_force[2054] <= 8'h64;
  filter_in_data_log_force[2055] <= 8'ha6;
  filter_in_data_log_force[2056] <= 8'h4f;
  filter_in_data_log_force[2057] <= 8'hbc;
  filter_in_data_log_force[2058] <= 8'h38;
  filter_in_data_log_force[2059] <= 8'hd4;
  filter_in_data_log_force[2060] <= 8'h1f;
  filter_in_data_log_force[2061] <= 8'hed;
  filter_in_data_log_force[2062] <= 8'h07;
  filter_in_data_log_force[2063] <= 8'h05;
  filter_in_data_log_force[2064] <= 8'hf0;
  filter_in_data_log_force[2065] <= 8'h1b;
  filter_in_data_log_force[2066] <= 8'hdb;
  filter_in_data_log_force[2067] <= 8'h2e;
  filter_in_data_log_force[2068] <= 8'hc9;
  filter_in_data_log_force[2069] <= 8'h40;
  filter_in_data_log_force[2070] <= 8'hb9;
  filter_in_data_log_force[2071] <= 8'h4e;
  filter_in_data_log_force[2072] <= 8'hab;
  filter_in_data_log_force[2073] <= 8'h00;
  filter_in_data_log_force[2074] <= 8'h00;
  filter_in_data_log_force[2075] <= 8'h00;
  filter_in_data_log_force[2076] <= 8'h00;
  filter_in_data_log_force[2077] <= 8'h00;
  filter_in_data_log_force[2078] <= 8'hc0;
  filter_in_data_log_force[2079] <= 8'hfa;
  filter_in_data_log_force[2080] <= 8'he6;
  filter_in_data_log_force[2081] <= 8'h19;
  filter_in_data_log_force[2082] <= 8'h4d;
  filter_in_data_log_force[2083] <= 8'h9b;
  filter_in_data_log_force[2084] <= 8'h52;
  filter_in_data_log_force[2085] <= 8'h57;
  filter_in_data_log_force[2086] <= 8'hdb;
  filter_in_data_log_force[2087] <= 8'hee;
  filter_in_data_log_force[2088] <= 8'h12;
  filter_in_data_log_force[2089] <= 8'h33;
  filter_in_data_log_force[2090] <= 8'h3e;
  filter_in_data_log_force[2091] <= 8'h42;
  filter_in_data_log_force[2092] <= 8'he4;
  filter_in_data_log_force[2093] <= 8'hee;
  filter_in_data_log_force[2094] <= 8'h75;
  filter_in_data_log_force[2095] <= 8'h13;
  filter_in_data_log_force[2096] <= 8'h5a;
  filter_in_data_log_force[2097] <= 8'hc7;
  filter_in_data_log_force[2098] <= 8'h1f;
  filter_in_data_log_force[2099] <= 8'h17;
  filter_in_data_log_force[2100] <= 8'h77;
  filter_in_data_log_force[2101] <= 8'h96;
  filter_in_data_log_force[2102] <= 8'h00;
  filter_in_data_log_force[2103] <= 8'h06;
  filter_in_data_log_force[2104] <= 8'h97;
  filter_in_data_log_force[2105] <= 8'h68;
  filter_in_data_log_force[2106] <= 8'h62;
  filter_in_data_log_force[2107] <= 8'hf0;
  filter_in_data_log_force[2108] <= 8'h48;
  filter_in_data_log_force[2109] <= 8'ha6;
  filter_in_data_log_force[2110] <= 8'h1f;
  filter_in_data_log_force[2111] <= 8'hc3;
  filter_in_data_log_force[2112] <= 8'hf2;
  filter_in_data_log_force[2113] <= 8'h58;
  filter_in_data_log_force[2114] <= 8'hb2;
  filter_in_data_log_force[2115] <= 8'hce;
  filter_in_data_log_force[2116] <= 8'hfc;
  filter_in_data_log_force[2117] <= 8'hd6;
  filter_in_data_log_force[2118] <= 8'h4c;
  filter_in_data_log_force[2119] <= 8'h7d;
  filter_in_data_log_force[2120] <= 8'ha9;
  filter_in_data_log_force[2121] <= 8'hbd;
  filter_in_data_log_force[2122] <= 8'h34;
  filter_in_data_log_force[2123] <= 8'he0;
  filter_in_data_log_force[2124] <= 8'h79;
  filter_in_data_log_force[2125] <= 8'h79;
  filter_in_data_log_force[2126] <= 8'h25;
  filter_in_data_log_force[2127] <= 8'h5c;
  filter_in_data_log_force[2128] <= 8'he7;
  filter_in_data_log_force[2129] <= 8'h22;
  filter_in_data_log_force[2130] <= 8'h7c;
  filter_in_data_log_force[2131] <= 8'h0f;
  filter_in_data_log_force[2132] <= 8'h6f;
  filter_in_data_log_force[2133] <= 8'h38;
  filter_in_data_log_force[2134] <= 8'hfc;
  filter_in_data_log_force[2135] <= 8'h24;
  filter_in_data_log_force[2136] <= 8'h63;
  filter_in_data_log_force[2137] <= 8'hb3;
  filter_in_data_log_force[2138] <= 8'he5;
  filter_in_data_log_force[2139] <= 8'h7e;
  filter_in_data_log_force[2140] <= 8'he7;
  filter_in_data_log_force[2141] <= 8'h29;
  filter_in_data_log_force[2142] <= 8'h67;
  filter_in_data_log_force[2143] <= 8'h7f;
  filter_in_data_log_force[2144] <= 8'h27;
  filter_in_data_log_force[2145] <= 8'h9c;
  filter_in_data_log_force[2146] <= 8'h89;
  filter_in_data_log_force[2147] <= 8'h1e;
  filter_in_data_log_force[2148] <= 8'h11;
  filter_in_data_log_force[2149] <= 8'h76;
  filter_in_data_log_force[2150] <= 8'h3f;
  filter_in_data_log_force[2151] <= 8'h2a;
  filter_in_data_log_force[2152] <= 8'h06;
  filter_in_data_log_force[2153] <= 8'hc3;
  filter_in_data_log_force[2154] <= 8'h76;
  filter_in_data_log_force[2155] <= 8'h0a;
  filter_in_data_log_force[2156] <= 8'h88;
  filter_in_data_log_force[2157] <= 8'h32;
  filter_in_data_log_force[2158] <= 8'h05;
  filter_in_data_log_force[2159] <= 8'h8f;
  filter_in_data_log_force[2160] <= 8'h64;
  filter_in_data_log_force[2161] <= 8'hd5;
  filter_in_data_log_force[2162] <= 8'hbb;
  filter_in_data_log_force[2163] <= 8'h9d;
  filter_in_data_log_force[2164] <= 8'hd0;
  filter_in_data_log_force[2165] <= 8'hba;
  filter_in_data_log_force[2166] <= 8'h27;
  filter_in_data_log_force[2167] <= 8'h91;
  filter_in_data_log_force[2168] <= 8'hc7;
  filter_in_data_log_force[2169] <= 8'hc8;
  filter_in_data_log_force[2170] <= 8'h61;
  filter_in_data_log_force[2171] <= 8'hf2;
  filter_in_data_log_force[2172] <= 8'h42;
  filter_in_data_log_force[2173] <= 8'h1a;
  filter_in_data_log_force[2174] <= 8'h49;
  filter_in_data_log_force[2175] <= 8'h9d;
  filter_in_data_log_force[2176] <= 8'h7b;
  filter_in_data_log_force[2177] <= 8'h59;
  filter_in_data_log_force[2178] <= 8'h8d;
  filter_in_data_log_force[2179] <= 8'hf7;
  filter_in_data_log_force[2180] <= 8'hd3;
  filter_in_data_log_force[2181] <= 8'h21;
  filter_in_data_log_force[2182] <= 8'hbb;
  filter_in_data_log_force[2183] <= 8'h14;
  filter_in_data_log_force[2184] <= 8'h1a;
  filter_in_data_log_force[2185] <= 8'h1a;
  filter_in_data_log_force[2186] <= 8'hf3;
  filter_in_data_log_force[2187] <= 8'h89;
  filter_in_data_log_force[2188] <= 8'h04;
  filter_in_data_log_force[2189] <= 8'he8;
  filter_in_data_log_force[2190] <= 8'h9c;
  filter_in_data_log_force[2191] <= 8'hf6;
  filter_in_data_log_force[2192] <= 8'hf3;
  filter_in_data_log_force[2193] <= 8'h0d;
  filter_in_data_log_force[2194] <= 8'h4e;
  filter_in_data_log_force[2195] <= 8'h33;
  filter_in_data_log_force[2196] <= 8'h5f;
  filter_in_data_log_force[2197] <= 8'h8d;
  filter_in_data_log_force[2198] <= 8'hb8;
  filter_in_data_log_force[2199] <= 8'hf6;
  filter_in_data_log_force[2200] <= 8'h75;
  filter_in_data_log_force[2201] <= 8'h4a;
  filter_in_data_log_force[2202] <= 8'hf4;
  filter_in_data_log_force[2203] <= 8'hd5;
  filter_in_data_log_force[2204] <= 8'h8f;
  filter_in_data_log_force[2205] <= 8'h3e;
  filter_in_data_log_force[2206] <= 8'h02;
  filter_in_data_log_force[2207] <= 8'hb3;
  filter_in_data_log_force[2208] <= 8'hed;
  filter_in_data_log_force[2209] <= 8'hab;
  filter_in_data_log_force[2210] <= 8'h40;
  filter_in_data_log_force[2211] <= 8'hde;
  filter_in_data_log_force[2212] <= 8'h71;
  filter_in_data_log_force[2213] <= 8'h84;
  filter_in_data_log_force[2214] <= 8'h54;
  filter_in_data_log_force[2215] <= 8'h20;
  filter_in_data_log_force[2216] <= 8'h0a;
  filter_in_data_log_force[2217] <= 8'h27;
  filter_in_data_log_force[2218] <= 8'h3a;
  filter_in_data_log_force[2219] <= 8'h98;
  filter_in_data_log_force[2220] <= 8'h61;
  filter_in_data_log_force[2221] <= 8'h84;
  filter_in_data_log_force[2222] <= 8'hcb;
  filter_in_data_log_force[2223] <= 8'hae;
  filter_in_data_log_force[2224] <= 8'h6d;
  filter_in_data_log_force[2225] <= 8'h91;
  filter_in_data_log_force[2226] <= 8'h15;
  filter_in_data_log_force[2227] <= 8'h23;
  filter_in_data_log_force[2228] <= 8'h27;
  filter_in_data_log_force[2229] <= 8'h5d;
  filter_in_data_log_force[2230] <= 8'h8e;
  filter_in_data_log_force[2231] <= 8'h51;
  filter_in_data_log_force[2232] <= 8'h07;
  filter_in_data_log_force[2233] <= 8'h32;
  filter_in_data_log_force[2234] <= 8'hb6;
  filter_in_data_log_force[2235] <= 8'h0b;
  filter_in_data_log_force[2236] <= 8'h34;
  filter_in_data_log_force[2237] <= 8'h75;
  filter_in_data_log_force[2238] <= 8'hf2;
  filter_in_data_log_force[2239] <= 8'h96;
  filter_in_data_log_force[2240] <= 8'h8f;
  filter_in_data_log_force[2241] <= 8'h21;
  filter_in_data_log_force[2242] <= 8'h4c;
  filter_in_data_log_force[2243] <= 8'h31;
  filter_in_data_log_force[2244] <= 8'hd8;
  filter_in_data_log_force[2245] <= 8'h72;
  filter_in_data_log_force[2246] <= 8'h05;
  filter_in_data_log_force[2247] <= 8'h74;
  filter_in_data_log_force[2248] <= 8'h93;
  filter_in_data_log_force[2249] <= 8'hb5;
  filter_in_data_log_force[2250] <= 8'h46;
  filter_in_data_log_force[2251] <= 8'h6a;
  filter_in_data_log_force[2252] <= 8'h48;
  filter_in_data_log_force[2253] <= 8'hcc;
  filter_in_data_log_force[2254] <= 8'ha7;
  filter_in_data_log_force[2255] <= 8'h59;
  filter_in_data_log_force[2256] <= 8'h49;
  filter_in_data_log_force[2257] <= 8'hc5;
  filter_in_data_log_force[2258] <= 8'hba;
  filter_in_data_log_force[2259] <= 8'hd2;
  filter_in_data_log_force[2260] <= 8'h54;
  filter_in_data_log_force[2261] <= 8'h52;
  filter_in_data_log_force[2262] <= 8'h12;
  filter_in_data_log_force[2263] <= 8'h12;
  filter_in_data_log_force[2264] <= 8'hc9;
  filter_in_data_log_force[2265] <= 8'h33;
  filter_in_data_log_force[2266] <= 8'h4c;
  filter_in_data_log_force[2267] <= 8'hf1;
  filter_in_data_log_force[2268] <= 8'hf2;
  filter_in_data_log_force[2269] <= 8'hf7;
  filter_in_data_log_force[2270] <= 8'hc7;
  filter_in_data_log_force[2271] <= 8'h2d;
  filter_in_data_log_force[2272] <= 8'h67;
  filter_in_data_log_force[2273] <= 8'h69;
  filter_in_data_log_force[2274] <= 8'h3f;
  filter_in_data_log_force[2275] <= 8'hc3;
  filter_in_data_log_force[2276] <= 8'h31;
  filter_in_data_log_force[2277] <= 8'ha2;
  filter_in_data_log_force[2278] <= 8'ha0;
  filter_in_data_log_force[2279] <= 8'hb1;
  filter_in_data_log_force[2280] <= 8'ha5;
  filter_in_data_log_force[2281] <= 8'h16;
  filter_in_data_log_force[2282] <= 8'h93;
  filter_in_data_log_force[2283] <= 8'h53;
  filter_in_data_log_force[2284] <= 8'h39;
  filter_in_data_log_force[2285] <= 8'h6d;
  filter_in_data_log_force[2286] <= 8'hfe;
  filter_in_data_log_force[2287] <= 8'h28;
  filter_in_data_log_force[2288] <= 8'h64;
  filter_in_data_log_force[2289] <= 8'h0a;
  filter_in_data_log_force[2290] <= 8'hc8;
  filter_in_data_log_force[2291] <= 8'h7a;
  filter_in_data_log_force[2292] <= 8'h89;
  filter_in_data_log_force[2293] <= 8'hd4;
  filter_in_data_log_force[2294] <= 8'h79;
  filter_in_data_log_force[2295] <= 8'hdd;
  filter_in_data_log_force[2296] <= 8'hcf;
  filter_in_data_log_force[2297] <= 8'h9f;
  filter_in_data_log_force[2298] <= 8'h6a;
  filter_in_data_log_force[2299] <= 8'ha3;
  filter_in_data_log_force[2300] <= 8'hd5;
  filter_in_data_log_force[2301] <= 8'h66;
  filter_in_data_log_force[2302] <= 8'h00;
  filter_in_data_log_force[2303] <= 8'h1e;
  filter_in_data_log_force[2304] <= 8'h15;
  filter_in_data_log_force[2305] <= 8'h33;
  filter_in_data_log_force[2306] <= 8'h88;
  filter_in_data_log_force[2307] <= 8'h07;
  filter_in_data_log_force[2308] <= 8'h88;
  filter_in_data_log_force[2309] <= 8'h54;
  filter_in_data_log_force[2310] <= 8'hd7;
  filter_in_data_log_force[2311] <= 8'h59;
  filter_in_data_log_force[2312] <= 8'hbf;
  filter_in_data_log_force[2313] <= 8'h15;
  filter_in_data_log_force[2314] <= 8'h70;
  filter_in_data_log_force[2315] <= 8'h8c;
  filter_in_data_log_force[2316] <= 8'h8e;
  filter_in_data_log_force[2317] <= 8'h85;
  filter_in_data_log_force[2318] <= 8'h2e;
  filter_in_data_log_force[2319] <= 8'h19;
  filter_in_data_log_force[2320] <= 8'h9d;
  filter_in_data_log_force[2321] <= 8'h4c;
  filter_in_data_log_force[2322] <= 8'h1e;
  filter_in_data_log_force[2323] <= 8'h92;
  filter_in_data_log_force[2324] <= 8'h92;
  filter_in_data_log_force[2325] <= 8'ha3;
  filter_in_data_log_force[2326] <= 8'h4a;
  filter_in_data_log_force[2327] <= 8'h98;
  filter_in_data_log_force[2328] <= 8'hbd;
  filter_in_data_log_force[2329] <= 8'hbe;
  filter_in_data_log_force[2330] <= 8'h9b;
  filter_in_data_log_force[2331] <= 8'h5c;
  filter_in_data_log_force[2332] <= 8'h33;
  filter_in_data_log_force[2333] <= 8'h3c;
  filter_in_data_log_force[2334] <= 8'h27;
  filter_in_data_log_force[2335] <= 8'h04;
  filter_in_data_log_force[2336] <= 8'hd4;
  filter_in_data_log_force[2337] <= 8'h29;
  filter_in_data_log_force[2338] <= 8'h9e;
  filter_in_data_log_force[2339] <= 8'ha6;
  filter_in_data_log_force[2340] <= 8'h85;
  filter_in_data_log_force[2341] <= 8'h77;
  filter_in_data_log_force[2342] <= 8'h78;
  filter_in_data_log_force[2343] <= 8'ha0;
  filter_in_data_log_force[2344] <= 8'hf8;
  filter_in_data_log_force[2345] <= 8'h28;
  filter_in_data_log_force[2346] <= 8'hca;
  filter_in_data_log_force[2347] <= 8'h41;
  filter_in_data_log_force[2348] <= 8'h0f;
  filter_in_data_log_force[2349] <= 8'hee;
  filter_in_data_log_force[2350] <= 8'hc4;
  filter_in_data_log_force[2351] <= 8'h41;
  filter_in_data_log_force[2352] <= 8'h66;
  filter_in_data_log_force[2353] <= 8'h3a;
  filter_in_data_log_force[2354] <= 8'he8;
  filter_in_data_log_force[2355] <= 8'h70;
  filter_in_data_log_force[2356] <= 8'hc1;
  filter_in_data_log_force[2357] <= 8'h08;
  filter_in_data_log_force[2358] <= 8'h74;
  filter_in_data_log_force[2359] <= 8'hc5;
  filter_in_data_log_force[2360] <= 8'hc0;
  filter_in_data_log_force[2361] <= 8'h6d;
  filter_in_data_log_force[2362] <= 8'h92;
  filter_in_data_log_force[2363] <= 8'hcd;
  filter_in_data_log_force[2364] <= 8'h17;
  filter_in_data_log_force[2365] <= 8'hb4;
  filter_in_data_log_force[2366] <= 8'h23;
  filter_in_data_log_force[2367] <= 8'h4c;
  filter_in_data_log_force[2368] <= 8'h00;
  filter_in_data_log_force[2369] <= 8'h27;
  filter_in_data_log_force[2370] <= 8'h4c;
  filter_in_data_log_force[2371] <= 8'hbc;
  filter_in_data_log_force[2372] <= 8'h1a;
  filter_in_data_log_force[2373] <= 8'h9d;
  filter_in_data_log_force[2374] <= 8'h04;
  filter_in_data_log_force[2375] <= 8'h56;
  filter_in_data_log_force[2376] <= 8'h6c;
  filter_in_data_log_force[2377] <= 8'h00;
  filter_in_data_log_force[2378] <= 8'hc7;
  filter_in_data_log_force[2379] <= 8'h27;
  filter_in_data_log_force[2380] <= 8'h6b;
  filter_in_data_log_force[2381] <= 8'h03;
  filter_in_data_log_force[2382] <= 8'h79;
  filter_in_data_log_force[2383] <= 8'hb3;
  filter_in_data_log_force[2384] <= 8'h9c;
  filter_in_data_log_force[2385] <= 8'hcc;
  filter_in_data_log_force[2386] <= 8'he5;
  filter_in_data_log_force[2387] <= 8'hec;
  filter_in_data_log_force[2388] <= 8'hd0;
  filter_in_data_log_force[2389] <= 8'h32;
  filter_in_data_log_force[2390] <= 8'h98;
  filter_in_data_log_force[2391] <= 8'he7;
  filter_in_data_log_force[2392] <= 8'hcc;
  filter_in_data_log_force[2393] <= 8'hce;
  filter_in_data_log_force[2394] <= 8'h9b;
  filter_in_data_log_force[2395] <= 8'h18;
  filter_in_data_log_force[2396] <= 8'hc8;
  filter_in_data_log_force[2397] <= 8'ha8;
  filter_in_data_log_force[2398] <= 8'h80;
  filter_in_data_log_force[2399] <= 8'hc9;
  filter_in_data_log_force[2400] <= 8'h0d;
  filter_in_data_log_force[2401] <= 8'h5f;
  filter_in_data_log_force[2402] <= 8'h8b;
  filter_in_data_log_force[2403] <= 8'h68;
  filter_in_data_log_force[2404] <= 8'ha2;
  filter_in_data_log_force[2405] <= 8'h55;
  filter_in_data_log_force[2406] <= 8'h4d;
  filter_in_data_log_force[2407] <= 8'h6b;
  filter_in_data_log_force[2408] <= 8'ha3;
  filter_in_data_log_force[2409] <= 8'h01;
  filter_in_data_log_force[2410] <= 8'he8;
  filter_in_data_log_force[2411] <= 8'hac;
  filter_in_data_log_force[2412] <= 8'h13;
  filter_in_data_log_force[2413] <= 8'h1b;
  filter_in_data_log_force[2414] <= 8'hb7;
  filter_in_data_log_force[2415] <= 8'h05;
  filter_in_data_log_force[2416] <= 8'h7d;
  filter_in_data_log_force[2417] <= 8'hfd;
  filter_in_data_log_force[2418] <= 8'h32;
  filter_in_data_log_force[2419] <= 8'he9;
  filter_in_data_log_force[2420] <= 8'h89;
  filter_in_data_log_force[2421] <= 8'hcb;
  filter_in_data_log_force[2422] <= 8'h4d;
  filter_in_data_log_force[2423] <= 8'hd9;
  filter_in_data_log_force[2424] <= 8'h95;
  filter_in_data_log_force[2425] <= 8'h03;
  filter_in_data_log_force[2426] <= 8'hde;
  filter_in_data_log_force[2427] <= 8'h3d;
  filter_in_data_log_force[2428] <= 8'h06;
  filter_in_data_log_force[2429] <= 8'h4e;
  filter_in_data_log_force[2430] <= 8'h51;
  filter_in_data_log_force[2431] <= 8'hb1;
  filter_in_data_log_force[2432] <= 8'ha0;
  filter_in_data_log_force[2433] <= 8'h52;
  filter_in_data_log_force[2434] <= 8'h23;
  filter_in_data_log_force[2435] <= 8'h84;
  filter_in_data_log_force[2436] <= 8'h65;
  filter_in_data_log_force[2437] <= 8'h04;
  filter_in_data_log_force[2438] <= 8'h0b;
  filter_in_data_log_force[2439] <= 8'h1b;
  filter_in_data_log_force[2440] <= 8'h43;
  filter_in_data_log_force[2441] <= 8'h5b;
  filter_in_data_log_force[2442] <= 8'he2;
  filter_in_data_log_force[2443] <= 8'h96;
  filter_in_data_log_force[2444] <= 8'h3c;
  filter_in_data_log_force[2445] <= 8'hd5;
  filter_in_data_log_force[2446] <= 8'h57;
  filter_in_data_log_force[2447] <= 8'hdf;
  filter_in_data_log_force[2448] <= 8'h54;
  filter_in_data_log_force[2449] <= 8'had;
  filter_in_data_log_force[2450] <= 8'ha1;
  filter_in_data_log_force[2451] <= 8'h61;
  filter_in_data_log_force[2452] <= 8'h8b;
  filter_in_data_log_force[2453] <= 8'h30;
  filter_in_data_log_force[2454] <= 8'h3c;
  filter_in_data_log_force[2455] <= 8'hf0;
  filter_in_data_log_force[2456] <= 8'he1;
  filter_in_data_log_force[2457] <= 8'h7b;
  filter_in_data_log_force[2458] <= 8'he6;
  filter_in_data_log_force[2459] <= 8'hf1;
  filter_in_data_log_force[2460] <= 8'ha8;
  filter_in_data_log_force[2461] <= 8'hd3;
  filter_in_data_log_force[2462] <= 8'hd0;
  filter_in_data_log_force[2463] <= 8'h65;
  filter_in_data_log_force[2464] <= 8'hbf;
  filter_in_data_log_force[2465] <= 8'hd0;
  filter_in_data_log_force[2466] <= 8'he9;
  filter_in_data_log_force[2467] <= 8'h35;
  filter_in_data_log_force[2468] <= 8'ha5;
  filter_in_data_log_force[2469] <= 8'h5f;
  filter_in_data_log_force[2470] <= 8'h95;
  filter_in_data_log_force[2471] <= 8'hf6;
  filter_in_data_log_force[2472] <= 8'h88;
  filter_in_data_log_force[2473] <= 8'h41;
  filter_in_data_log_force[2474] <= 8'h33;
  filter_in_data_log_force[2475] <= 8'hb7;
  filter_in_data_log_force[2476] <= 8'h2e;
  filter_in_data_log_force[2477] <= 8'h0f;
  filter_in_data_log_force[2478] <= 8'h5a;
  filter_in_data_log_force[2479] <= 8'h0f;
  filter_in_data_log_force[2480] <= 8'h67;
  filter_in_data_log_force[2481] <= 8'heb;
  filter_in_data_log_force[2482] <= 8'hdc;
  filter_in_data_log_force[2483] <= 8'hfd;
  filter_in_data_log_force[2484] <= 8'hc2;
  filter_in_data_log_force[2485] <= 8'h6e;
  filter_in_data_log_force[2486] <= 8'hf7;
  filter_in_data_log_force[2487] <= 8'hc1;
  filter_in_data_log_force[2488] <= 8'hee;
  filter_in_data_log_force[2489] <= 8'h34;
  filter_in_data_log_force[2490] <= 8'he7;
  filter_in_data_log_force[2491] <= 8'haf;
  filter_in_data_log_force[2492] <= 8'h5b;
  filter_in_data_log_force[2493] <= 8'h16;
  filter_in_data_log_force[2494] <= 8'he0;
  filter_in_data_log_force[2495] <= 8'hb9;
  filter_in_data_log_force[2496] <= 8'hb8;
  filter_in_data_log_force[2497] <= 8'h06;
  filter_in_data_log_force[2498] <= 8'hef;
  filter_in_data_log_force[2499] <= 8'h3e;
  filter_in_data_log_force[2500] <= 8'h92;
  filter_in_data_log_force[2501] <= 8'h59;
  filter_in_data_log_force[2502] <= 8'h2e;
  filter_in_data_log_force[2503] <= 8'ha3;
  filter_in_data_log_force[2504] <= 8'h5c;
  filter_in_data_log_force[2505] <= 8'hb3;
  filter_in_data_log_force[2506] <= 8'h1b;
  filter_in_data_log_force[2507] <= 8'h0b;
  filter_in_data_log_force[2508] <= 8'haa;
  filter_in_data_log_force[2509] <= 8'h81;
  filter_in_data_log_force[2510] <= 8'h46;
  filter_in_data_log_force[2511] <= 8'h44;
  filter_in_data_log_force[2512] <= 8'hec;
  filter_in_data_log_force[2513] <= 8'h8f;
  filter_in_data_log_force[2514] <= 8'h16;
  filter_in_data_log_force[2515] <= 8'had;
  filter_in_data_log_force[2516] <= 8'h3b;
  filter_in_data_log_force[2517] <= 8'h09;
  filter_in_data_log_force[2518] <= 8'hc1;
  filter_in_data_log_force[2519] <= 8'h6b;
  filter_in_data_log_force[2520] <= 8'h42;
  filter_in_data_log_force[2521] <= 8'h63;
  filter_in_data_log_force[2522] <= 8'h92;
  filter_in_data_log_force[2523] <= 8'haf;
  filter_in_data_log_force[2524] <= 8'h3d;
  filter_in_data_log_force[2525] <= 8'h32;
  filter_in_data_log_force[2526] <= 8'h47;
  filter_in_data_log_force[2527] <= 8'h00;
  filter_in_data_log_force[2528] <= 8'hed;
  filter_in_data_log_force[2529] <= 8'h1c;
  filter_in_data_log_force[2530] <= 8'h5b;
  filter_in_data_log_force[2531] <= 8'h2c;
  filter_in_data_log_force[2532] <= 8'h06;
  filter_in_data_log_force[2533] <= 8'hcc;
  filter_in_data_log_force[2534] <= 8'h34;
  filter_in_data_log_force[2535] <= 8'he2;
  filter_in_data_log_force[2536] <= 8'h11;
  filter_in_data_log_force[2537] <= 8'h63;
  filter_in_data_log_force[2538] <= 8'h58;
  filter_in_data_log_force[2539] <= 8'h66;
  filter_in_data_log_force[2540] <= 8'h70;
  filter_in_data_log_force[2541] <= 8'h51;
  filter_in_data_log_force[2542] <= 8'h80;
  filter_in_data_log_force[2543] <= 8'h81;
  filter_in_data_log_force[2544] <= 8'h96;
  filter_in_data_log_force[2545] <= 8'hc3;
  filter_in_data_log_force[2546] <= 8'h86;
  filter_in_data_log_force[2547] <= 8'hed;
  filter_in_data_log_force[2548] <= 8'hd7;
  filter_in_data_log_force[2549] <= 8'h0b;
  filter_in_data_log_force[2550] <= 8'h6d;
  filter_in_data_log_force[2551] <= 8'hcc;
  filter_in_data_log_force[2552] <= 8'hd7;
  filter_in_data_log_force[2553] <= 8'h5c;
  filter_in_data_log_force[2554] <= 8'hd7;
  filter_in_data_log_force[2555] <= 8'ha3;
  filter_in_data_log_force[2556] <= 8'h02;
  filter_in_data_log_force[2557] <= 8'h5b;
  filter_in_data_log_force[2558] <= 8'he2;
  filter_in_data_log_force[2559] <= 8'h32;
  filter_in_data_log_force[2560] <= 8'h21;
  filter_in_data_log_force[2561] <= 8'hf3;
  filter_in_data_log_force[2562] <= 8'hf9;
  filter_in_data_log_force[2563] <= 8'h73;
  filter_in_data_log_force[2564] <= 8'h95;
  filter_in_data_log_force[2565] <= 8'hc8;
  filter_in_data_log_force[2566] <= 8'hf2;
  filter_in_data_log_force[2567] <= 8'h16;
  filter_in_data_log_force[2568] <= 8'h61;
  filter_in_data_log_force[2569] <= 8'hf8;
  filter_in_data_log_force[2570] <= 8'hf0;
  filter_in_data_log_force[2571] <= 8'h3f;
  filter_in_data_log_force[2572] <= 8'hf8;
  filter_in_data_log_force[2573] <= 8'h5c;
  filter_in_data_log_force[2574] <= 8'hf7;
  filter_in_data_log_force[2575] <= 8'h00;
  filter_in_data_log_force[2576] <= 8'hfd;
  filter_in_data_log_force[2577] <= 8'hbb;
  filter_in_data_log_force[2578] <= 8'h96;
  filter_in_data_log_force[2579] <= 8'h91;
  filter_in_data_log_force[2580] <= 8'h63;
  filter_in_data_log_force[2581] <= 8'hbc;
  filter_in_data_log_force[2582] <= 8'h5d;
  filter_in_data_log_force[2583] <= 8'h36;
  filter_in_data_log_force[2584] <= 8'h5f;
  filter_in_data_log_force[2585] <= 8'h70;
  filter_in_data_log_force[2586] <= 8'ha4;
  filter_in_data_log_force[2587] <= 8'he5;
  filter_in_data_log_force[2588] <= 8'h7b;
  filter_in_data_log_force[2589] <= 8'h25;
  filter_in_data_log_force[2590] <= 8'h65;
  filter_in_data_log_force[2591] <= 8'hfb;
  filter_in_data_log_force[2592] <= 8'h84;
  filter_in_data_log_force[2593] <= 8'h1f;
  filter_in_data_log_force[2594] <= 8'hbb;
  filter_in_data_log_force[2595] <= 8'h07;
  filter_in_data_log_force[2596] <= 8'h3a;
  filter_in_data_log_force[2597] <= 8'h1b;
  filter_in_data_log_force[2598] <= 8'h17;
  filter_in_data_log_force[2599] <= 8'hef;
  filter_in_data_log_force[2600] <= 8'hbf;
  filter_in_data_log_force[2601] <= 8'hee;
  filter_in_data_log_force[2602] <= 8'h83;
  filter_in_data_log_force[2603] <= 8'h1c;
  filter_in_data_log_force[2604] <= 8'h75;
  filter_in_data_log_force[2605] <= 8'h98;
  filter_in_data_log_force[2606] <= 8'h89;
  filter_in_data_log_force[2607] <= 8'h63;
  filter_in_data_log_force[2608] <= 8'hbf;
  filter_in_data_log_force[2609] <= 8'h82;
  filter_in_data_log_force[2610] <= 8'h51;
  filter_in_data_log_force[2611] <= 8'ha4;
  filter_in_data_log_force[2612] <= 8'h61;
  filter_in_data_log_force[2613] <= 8'h98;
  filter_in_data_log_force[2614] <= 8'hda;
  filter_in_data_log_force[2615] <= 8'h18;
  filter_in_data_log_force[2616] <= 8'h16;
  filter_in_data_log_force[2617] <= 8'h2b;
  filter_in_data_log_force[2618] <= 8'h26;
  filter_in_data_log_force[2619] <= 8'hef;
  filter_in_data_log_force[2620] <= 8'ha4;
  filter_in_data_log_force[2621] <= 8'h40;
  filter_in_data_log_force[2622] <= 8'hbe;
  filter_in_data_log_force[2623] <= 8'h27;
  filter_in_data_log_force[2624] <= 8'h5b;
  filter_in_data_log_force[2625] <= 8'h96;
  filter_in_data_log_force[2626] <= 8'h79;
  filter_in_data_log_force[2627] <= 8'h88;
  filter_in_data_log_force[2628] <= 8'h56;
  filter_in_data_log_force[2629] <= 8'h56;
  filter_in_data_log_force[2630] <= 8'h8d;
  filter_in_data_log_force[2631] <= 8'h0c;
  filter_in_data_log_force[2632] <= 8'h71;
  filter_in_data_log_force[2633] <= 8'hd2;
  filter_in_data_log_force[2634] <= 8'h4e;
  filter_in_data_log_force[2635] <= 8'h1a;
  filter_in_data_log_force[2636] <= 8'h4a;
  filter_in_data_log_force[2637] <= 8'h4d;
  filter_in_data_log_force[2638] <= 8'h8d;
  filter_in_data_log_force[2639] <= 8'hc8;
  filter_in_data_log_force[2640] <= 8'h27;
  filter_in_data_log_force[2641] <= 8'hfd;
  filter_in_data_log_force[2642] <= 8'h79;
  filter_in_data_log_force[2643] <= 8'h40;
  filter_in_data_log_force[2644] <= 8'h11;
  filter_in_data_log_force[2645] <= 8'hcd;
  filter_in_data_log_force[2646] <= 8'hc2;
  filter_in_data_log_force[2647] <= 8'h63;
  filter_in_data_log_force[2648] <= 8'hf2;
  filter_in_data_log_force[2649] <= 8'h51;
  filter_in_data_log_force[2650] <= 8'h99;
  filter_in_data_log_force[2651] <= 8'h5c;
  filter_in_data_log_force[2652] <= 8'h87;
  filter_in_data_log_force[2653] <= 8'h66;
  filter_in_data_log_force[2654] <= 8'h66;
  filter_in_data_log_force[2655] <= 8'h06;
  filter_in_data_log_force[2656] <= 8'h9f;
  filter_in_data_log_force[2657] <= 8'hae;
  filter_in_data_log_force[2658] <= 8'h35;
  filter_in_data_log_force[2659] <= 8'h55;
  filter_in_data_log_force[2660] <= 8'h89;
  filter_in_data_log_force[2661] <= 8'h42;
  filter_in_data_log_force[2662] <= 8'h75;
  filter_in_data_log_force[2663] <= 8'hd8;
  filter_in_data_log_force[2664] <= 8'h23;
  filter_in_data_log_force[2665] <= 8'hd8;
  filter_in_data_log_force[2666] <= 8'hb7;
  filter_in_data_log_force[2667] <= 8'h49;
  filter_in_data_log_force[2668] <= 8'h39;
  filter_in_data_log_force[2669] <= 8'hc7;
  filter_in_data_log_force[2670] <= 8'h15;
  filter_in_data_log_force[2671] <= 8'hec;
  filter_in_data_log_force[2672] <= 8'h98;
  filter_in_data_log_force[2673] <= 8'h86;
  filter_in_data_log_force[2674] <= 8'hfe;
  filter_in_data_log_force[2675] <= 8'hc7;
  filter_in_data_log_force[2676] <= 8'hd7;
  filter_in_data_log_force[2677] <= 8'hca;
  filter_in_data_log_force[2678] <= 8'hac;
  filter_in_data_log_force[2679] <= 8'he6;
  filter_in_data_log_force[2680] <= 8'h33;
  filter_in_data_log_force[2681] <= 8'hb4;
  filter_in_data_log_force[2682] <= 8'h2b;
  filter_in_data_log_force[2683] <= 8'hf1;
  filter_in_data_log_force[2684] <= 8'hef;
  filter_in_data_log_force[2685] <= 8'had;
  filter_in_data_log_force[2686] <= 8'hb1;
  filter_in_data_log_force[2687] <= 8'h1e;
  filter_in_data_log_force[2688] <= 8'hc5;
  filter_in_data_log_force[2689] <= 8'h0f;
  filter_in_data_log_force[2690] <= 8'h72;
  filter_in_data_log_force[2691] <= 8'h37;
  filter_in_data_log_force[2692] <= 8'h2e;
  filter_in_data_log_force[2693] <= 8'h76;
  filter_in_data_log_force[2694] <= 8'h46;
  filter_in_data_log_force[2695] <= 8'h1c;
  filter_in_data_log_force[2696] <= 8'h73;
  filter_in_data_log_force[2697] <= 8'h8f;
  filter_in_data_log_force[2698] <= 8'hc5;
  filter_in_data_log_force[2699] <= 8'h7d;
  filter_in_data_log_force[2700] <= 8'h46;
  filter_in_data_log_force[2701] <= 8'hfa;
  filter_in_data_log_force[2702] <= 8'h2e;
  filter_in_data_log_force[2703] <= 8'heb;
  filter_in_data_log_force[2704] <= 8'he1;
  filter_in_data_log_force[2705] <= 8'hb7;
  filter_in_data_log_force[2706] <= 8'he2;
  filter_in_data_log_force[2707] <= 8'h88;
  filter_in_data_log_force[2708] <= 8'hf9;
  filter_in_data_log_force[2709] <= 8'hd5;
  filter_in_data_log_force[2710] <= 8'h7a;
  filter_in_data_log_force[2711] <= 8'h0e;
  filter_in_data_log_force[2712] <= 8'h59;
  filter_in_data_log_force[2713] <= 8'he8;
  filter_in_data_log_force[2714] <= 8'hf6;
  filter_in_data_log_force[2715] <= 8'h54;
  filter_in_data_log_force[2716] <= 8'h7e;
  filter_in_data_log_force[2717] <= 8'h06;
  filter_in_data_log_force[2718] <= 8'h6d;
  filter_in_data_log_force[2719] <= 8'h3d;
  filter_in_data_log_force[2720] <= 8'h11;
  filter_in_data_log_force[2721] <= 8'h78;
  filter_in_data_log_force[2722] <= 8'h53;
  filter_in_data_log_force[2723] <= 8'h76;
  filter_in_data_log_force[2724] <= 8'h25;
  filter_in_data_log_force[2725] <= 8'he1;
  filter_in_data_log_force[2726] <= 8'hfa;
  filter_in_data_log_force[2727] <= 8'h69;
  filter_in_data_log_force[2728] <= 8'h84;
  filter_in_data_log_force[2729] <= 8'ha8;
  filter_in_data_log_force[2730] <= 8'hf9;
  filter_in_data_log_force[2731] <= 8'h0b;
  filter_in_data_log_force[2732] <= 8'h8f;
  filter_in_data_log_force[2733] <= 8'h28;
  filter_in_data_log_force[2734] <= 8'h64;
  filter_in_data_log_force[2735] <= 8'h9c;
  filter_in_data_log_force[2736] <= 8'hf0;
  filter_in_data_log_force[2737] <= 8'hc8;
  filter_in_data_log_force[2738] <= 8'h7c;
  filter_in_data_log_force[2739] <= 8'h1c;
  filter_in_data_log_force[2740] <= 8'hc1;
  filter_in_data_log_force[2741] <= 8'ha2;
  filter_in_data_log_force[2742] <= 8'h0c;
  filter_in_data_log_force[2743] <= 8'h54;
  filter_in_data_log_force[2744] <= 8'h56;
  filter_in_data_log_force[2745] <= 8'h55;
  filter_in_data_log_force[2746] <= 8'hb4;
  filter_in_data_log_force[2747] <= 8'h0b;
  filter_in_data_log_force[2748] <= 8'h60;
  filter_in_data_log_force[2749] <= 8'h9f;
  filter_in_data_log_force[2750] <= 8'h5b;
  filter_in_data_log_force[2751] <= 8'h66;
  filter_in_data_log_force[2752] <= 8'hb8;
  filter_in_data_log_force[2753] <= 8'h94;
  filter_in_data_log_force[2754] <= 8'hf9;
  filter_in_data_log_force[2755] <= 8'h56;
  filter_in_data_log_force[2756] <= 8'hf8;
  filter_in_data_log_force[2757] <= 8'hea;
  filter_in_data_log_force[2758] <= 8'h01;
  filter_in_data_log_force[2759] <= 8'ha0;
  filter_in_data_log_force[2760] <= 8'ha2;
  filter_in_data_log_force[2761] <= 8'h5f;
  filter_in_data_log_force[2762] <= 8'h1a;
  filter_in_data_log_force[2763] <= 8'hc4;
  filter_in_data_log_force[2764] <= 8'h5d;
  filter_in_data_log_force[2765] <= 8'h8f;
  filter_in_data_log_force[2766] <= 8'hf5;
  filter_in_data_log_force[2767] <= 8'h39;
  filter_in_data_log_force[2768] <= 8'hd7;
  filter_in_data_log_force[2769] <= 8'he7;
  filter_in_data_log_force[2770] <= 8'h07;
  filter_in_data_log_force[2771] <= 8'h65;
  filter_in_data_log_force[2772] <= 8'h47;
  filter_in_data_log_force[2773] <= 8'h92;
  filter_in_data_log_force[2774] <= 8'hc7;
  filter_in_data_log_force[2775] <= 8'he1;
  filter_in_data_log_force[2776] <= 8'h5d;
  filter_in_data_log_force[2777] <= 8'hec;
  filter_in_data_log_force[2778] <= 8'hbd;
  filter_in_data_log_force[2779] <= 8'h19;
  filter_in_data_log_force[2780] <= 8'hfb;
  filter_in_data_log_force[2781] <= 8'h66;
  filter_in_data_log_force[2782] <= 8'h6f;
  filter_in_data_log_force[2783] <= 8'h51;
  filter_in_data_log_force[2784] <= 8'h35;
  filter_in_data_log_force[2785] <= 8'h3e;
  filter_in_data_log_force[2786] <= 8'h66;
  filter_in_data_log_force[2787] <= 8'h91;
  filter_in_data_log_force[2788] <= 8'hd6;
  filter_in_data_log_force[2789] <= 8'h81;
  filter_in_data_log_force[2790] <= 8'h54;
  filter_in_data_log_force[2791] <= 8'h02;
  filter_in_data_log_force[2792] <= 8'hde;
  filter_in_data_log_force[2793] <= 8'hba;
  filter_in_data_log_force[2794] <= 8'h09;
  filter_in_data_log_force[2795] <= 8'hca;
  filter_in_data_log_force[2796] <= 8'h92;
  filter_in_data_log_force[2797] <= 8'h96;
  filter_in_data_log_force[2798] <= 8'h91;
  filter_in_data_log_force[2799] <= 8'he9;
  filter_in_data_log_force[2800] <= 8'ha0;
  filter_in_data_log_force[2801] <= 8'hf1;
  filter_in_data_log_force[2802] <= 8'h66;
  filter_in_data_log_force[2803] <= 8'hdb;
  filter_in_data_log_force[2804] <= 8'h9f;
  filter_in_data_log_force[2805] <= 8'h12;
  filter_in_data_log_force[2806] <= 8'h60;
  filter_in_data_log_force[2807] <= 8'hd9;
  filter_in_data_log_force[2808] <= 8'h8b;
  filter_in_data_log_force[2809] <= 8'ha4;
  filter_in_data_log_force[2810] <= 8'h94;
  filter_in_data_log_force[2811] <= 8'h3e;
  filter_in_data_log_force[2812] <= 8'hf5;
  filter_in_data_log_force[2813] <= 8'h2b;
  filter_in_data_log_force[2814] <= 8'h33;
  filter_in_data_log_force[2815] <= 8'h12;
  filter_in_data_log_force[2816] <= 8'h21;
  filter_in_data_log_force[2817] <= 8'h61;
  filter_in_data_log_force[2818] <= 8'h2a;
  filter_in_data_log_force[2819] <= 8'h60;
  filter_in_data_log_force[2820] <= 8'hf8;
  filter_in_data_log_force[2821] <= 8'ha4;
  filter_in_data_log_force[2822] <= 8'h91;
  filter_in_data_log_force[2823] <= 8'h37;
  filter_in_data_log_force[2824] <= 8'hcf;
  filter_in_data_log_force[2825] <= 8'h2c;
  filter_in_data_log_force[2826] <= 8'h27;
  filter_in_data_log_force[2827] <= 8'h08;
  filter_in_data_log_force[2828] <= 8'h37;
  filter_in_data_log_force[2829] <= 8'h01;
  filter_in_data_log_force[2830] <= 8'hfd;
  filter_in_data_log_force[2831] <= 8'hff;
  filter_in_data_log_force[2832] <= 8'h70;
  filter_in_data_log_force[2833] <= 8'he4;
  filter_in_data_log_force[2834] <= 8'h9e;
  filter_in_data_log_force[2835] <= 8'hbe;
  filter_in_data_log_force[2836] <= 8'h2f;
  filter_in_data_log_force[2837] <= 8'h57;
  filter_in_data_log_force[2838] <= 8'h78;
  filter_in_data_log_force[2839] <= 8'hb7;
  filter_in_data_log_force[2840] <= 8'h43;
  filter_in_data_log_force[2841] <= 8'h16;
  filter_in_data_log_force[2842] <= 8'he7;
  filter_in_data_log_force[2843] <= 8'h03;
  filter_in_data_log_force[2844] <= 8'hff;
  filter_in_data_log_force[2845] <= 8'h27;
  filter_in_data_log_force[2846] <= 8'h3e;
  filter_in_data_log_force[2847] <= 8'hcd;
  filter_in_data_log_force[2848] <= 8'h97;
  filter_in_data_log_force[2849] <= 8'h53;
  filter_in_data_log_force[2850] <= 8'he4;
  filter_in_data_log_force[2851] <= 8'h46;
  filter_in_data_log_force[2852] <= 8'hae;
  filter_in_data_log_force[2853] <= 8'h9c;
  filter_in_data_log_force[2854] <= 8'h68;
  filter_in_data_log_force[2855] <= 8'h60;
  filter_in_data_log_force[2856] <= 8'h7f;
  filter_in_data_log_force[2857] <= 8'h5d;
  filter_in_data_log_force[2858] <= 8'h89;
  filter_in_data_log_force[2859] <= 8'h0b;
  filter_in_data_log_force[2860] <= 8'h7f;
  filter_in_data_log_force[2861] <= 8'h03;
  filter_in_data_log_force[2862] <= 8'h60;
  filter_in_data_log_force[2863] <= 8'h92;
  filter_in_data_log_force[2864] <= 8'h7d;
  filter_in_data_log_force[2865] <= 8'h6c;
  filter_in_data_log_force[2866] <= 8'h10;
  filter_in_data_log_force[2867] <= 8'hee;
  filter_in_data_log_force[2868] <= 8'hd6;
  filter_in_data_log_force[2869] <= 8'h39;
  filter_in_data_log_force[2870] <= 8'h83;
  filter_in_data_log_force[2871] <= 8'he0;
  filter_in_data_log_force[2872] <= 8'h6c;
  filter_in_data_log_force[2873] <= 8'h0c;
  filter_in_data_log_force[2874] <= 8'hf9;
  filter_in_data_log_force[2875] <= 8'hff;
  filter_in_data_log_force[2876] <= 8'hcf;
  filter_in_data_log_force[2877] <= 8'h73;
  filter_in_data_log_force[2878] <= 8'h7b;
  filter_in_data_log_force[2879] <= 8'h03;
  filter_in_data_log_force[2880] <= 8'h7e;
  filter_in_data_log_force[2881] <= 8'hf5;
  filter_in_data_log_force[2882] <= 8'hed;
  filter_in_data_log_force[2883] <= 8'hb7;
  filter_in_data_log_force[2884] <= 8'hb1;
  filter_in_data_log_force[2885] <= 8'h55;
  filter_in_data_log_force[2886] <= 8'h3a;
  filter_in_data_log_force[2887] <= 8'h08;
  filter_in_data_log_force[2888] <= 8'h54;
  filter_in_data_log_force[2889] <= 8'h03;
  filter_in_data_log_force[2890] <= 8'h0d;
  filter_in_data_log_force[2891] <= 8'hb7;
  filter_in_data_log_force[2892] <= 8'h16;
  filter_in_data_log_force[2893] <= 8'ha5;
  filter_in_data_log_force[2894] <= 8'h8d;
  filter_in_data_log_force[2895] <= 8'h2f;
  filter_in_data_log_force[2896] <= 8'h1c;
  filter_in_data_log_force[2897] <= 8'hb8;
  filter_in_data_log_force[2898] <= 8'he8;
  filter_in_data_log_force[2899] <= 8'h21;
  filter_in_data_log_force[2900] <= 8'h0e;
  filter_in_data_log_force[2901] <= 8'ha1;
  filter_in_data_log_force[2902] <= 8'hab;
  filter_in_data_log_force[2903] <= 8'h80;
  filter_in_data_log_force[2904] <= 8'heb;
  filter_in_data_log_force[2905] <= 8'hfd;
  filter_in_data_log_force[2906] <= 8'ha9;
  filter_in_data_log_force[2907] <= 8'h2b;
  filter_in_data_log_force[2908] <= 8'h85;
  filter_in_data_log_force[2909] <= 8'h9f;
  filter_in_data_log_force[2910] <= 8'h74;
  filter_in_data_log_force[2911] <= 8'h7a;
  filter_in_data_log_force[2912] <= 8'h88;
  filter_in_data_log_force[2913] <= 8'hfe;
  filter_in_data_log_force[2914] <= 8'h5d;
  filter_in_data_log_force[2915] <= 8'hbe;
  filter_in_data_log_force[2916] <= 8'h56;
  filter_in_data_log_force[2917] <= 8'h50;
  filter_in_data_log_force[2918] <= 8'h21;
  filter_in_data_log_force[2919] <= 8'h81;
  filter_in_data_log_force[2920] <= 8'he1;
  filter_in_data_log_force[2921] <= 8'h68;
  filter_in_data_log_force[2922] <= 8'h2e;
  filter_in_data_log_force[2923] <= 8'he1;
  filter_in_data_log_force[2924] <= 8'h22;
  filter_in_data_log_force[2925] <= 8'hbe;
  filter_in_data_log_force[2926] <= 8'h12;
  filter_in_data_log_force[2927] <= 8'h7b;
  filter_in_data_log_force[2928] <= 8'h5a;
  filter_in_data_log_force[2929] <= 8'hc9;
  filter_in_data_log_force[2930] <= 8'h2f;
  filter_in_data_log_force[2931] <= 8'hdc;
  filter_in_data_log_force[2932] <= 8'h7d;
  filter_in_data_log_force[2933] <= 8'h96;
  filter_in_data_log_force[2934] <= 8'hc0;
  filter_in_data_log_force[2935] <= 8'h50;
  filter_in_data_log_force[2936] <= 8'h96;
  filter_in_data_log_force[2937] <= 8'h08;
  filter_in_data_log_force[2938] <= 8'h4d;
  filter_in_data_log_force[2939] <= 8'h3d;
  filter_in_data_log_force[2940] <= 8'ha4;
  filter_in_data_log_force[2941] <= 8'hf0;
  filter_in_data_log_force[2942] <= 8'hda;
  filter_in_data_log_force[2943] <= 8'hfa;
  filter_in_data_log_force[2944] <= 8'h16;
  filter_in_data_log_force[2945] <= 8'ha5;
  filter_in_data_log_force[2946] <= 8'h68;
  filter_in_data_log_force[2947] <= 8'h24;
  filter_in_data_log_force[2948] <= 8'haa;
  filter_in_data_log_force[2949] <= 8'h11;
  filter_in_data_log_force[2950] <= 8'h6e;
  filter_in_data_log_force[2951] <= 8'h48;
  filter_in_data_log_force[2952] <= 8'h30;
  filter_in_data_log_force[2953] <= 8'hf7;
  filter_in_data_log_force[2954] <= 8'hc3;
  filter_in_data_log_force[2955] <= 8'h12;
  filter_in_data_log_force[2956] <= 8'hc0;
  filter_in_data_log_force[2957] <= 8'hd2;
  filter_in_data_log_force[2958] <= 8'h69;
  filter_in_data_log_force[2959] <= 8'h63;
  filter_in_data_log_force[2960] <= 8'h4b;
  filter_in_data_log_force[2961] <= 8'h6d;
  filter_in_data_log_force[2962] <= 8'hae;
  filter_in_data_log_force[2963] <= 8'h04;
  filter_in_data_log_force[2964] <= 8'h21;
  filter_in_data_log_force[2965] <= 8'h6a;
  filter_in_data_log_force[2966] <= 8'h2a;
  filter_in_data_log_force[2967] <= 8'he4;
  filter_in_data_log_force[2968] <= 8'h3d;
  filter_in_data_log_force[2969] <= 8'h51;
  filter_in_data_log_force[2970] <= 8'h1a;
  filter_in_data_log_force[2971] <= 8'h96;
  filter_in_data_log_force[2972] <= 8'h6c;
  filter_in_data_log_force[2973] <= 8'h8e;
  filter_in_data_log_force[2974] <= 8'h07;
  filter_in_data_log_force[2975] <= 8'h9e;
  filter_in_data_log_force[2976] <= 8'he1;
  filter_in_data_log_force[2977] <= 8'h50;
  filter_in_data_log_force[2978] <= 8'hbe;
  filter_in_data_log_force[2979] <= 8'h62;
  filter_in_data_log_force[2980] <= 8'h36;
  filter_in_data_log_force[2981] <= 8'he1;
  filter_in_data_log_force[2982] <= 8'hc0;
  filter_in_data_log_force[2983] <= 8'hc1;
  filter_in_data_log_force[2984] <= 8'h44;
  filter_in_data_log_force[2985] <= 8'h8d;
  filter_in_data_log_force[2986] <= 8'h2f;
  filter_in_data_log_force[2987] <= 8'h1f;
  filter_in_data_log_force[2988] <= 8'h3f;
  filter_in_data_log_force[2989] <= 8'h7a;
  filter_in_data_log_force[2990] <= 8'he2;
  filter_in_data_log_force[2991] <= 8'hc3;
  filter_in_data_log_force[2992] <= 8'h61;
  filter_in_data_log_force[2993] <= 8'h4e;
  filter_in_data_log_force[2994] <= 8'hf6;
  filter_in_data_log_force[2995] <= 8'h97;
  filter_in_data_log_force[2996] <= 8'h10;
  filter_in_data_log_force[2997] <= 8'hb0;
  filter_in_data_log_force[2998] <= 8'h08;
  filter_in_data_log_force[2999] <= 8'hdb;
  filter_in_data_log_force[3000] <= 8'hd1;
  filter_in_data_log_force[3001] <= 8'h3a;
  filter_in_data_log_force[3002] <= 8'h04;
  filter_in_data_log_force[3003] <= 8'h4a;
  filter_in_data_log_force[3004] <= 8'hb4;
  filter_in_data_log_force[3005] <= 8'h2e;
  filter_in_data_log_force[3006] <= 8'h8d;
  filter_in_data_log_force[3007] <= 8'h4d;
  filter_in_data_log_force[3008] <= 8'h2e;
  filter_in_data_log_force[3009] <= 8'h72;
  filter_in_data_log_force[3010] <= 8'h97;
  filter_in_data_log_force[3011] <= 8'h69;
  filter_in_data_log_force[3012] <= 8'h03;
  filter_in_data_log_force[3013] <= 8'h1d;
  filter_in_data_log_force[3014] <= 8'hd1;
  filter_in_data_log_force[3015] <= 8'h94;
  filter_in_data_log_force[3016] <= 8'h5a;
  filter_in_data_log_force[3017] <= 8'ha5;
  filter_in_data_log_force[3018] <= 8'hdf;
  filter_in_data_log_force[3019] <= 8'h1f;
  filter_in_data_log_force[3020] <= 8'h7f;
  filter_in_data_log_force[3021] <= 8'h04;
  filter_in_data_log_force[3022] <= 8'h7e;
  filter_in_data_log_force[3023] <= 8'hba;
  filter_in_data_log_force[3024] <= 8'he6;
  filter_in_data_log_force[3025] <= 8'h32;
  filter_in_data_log_force[3026] <= 8'h91;
  filter_in_data_log_force[3027] <= 8'h3f;
  filter_in_data_log_force[3028] <= 8'hec;
  filter_in_data_log_force[3029] <= 8'h50;
  filter_in_data_log_force[3030] <= 8'he1;
  filter_in_data_log_force[3031] <= 8'hd2;
  filter_in_data_log_force[3032] <= 8'h7c;
  filter_in_data_log_force[3033] <= 8'h38;
  filter_in_data_log_force[3034] <= 8'hea;
  filter_in_data_log_force[3035] <= 8'h99;
  filter_in_data_log_force[3036] <= 8'h3c;
  filter_in_data_log_force[3037] <= 8'h23;
  filter_in_data_log_force[3038] <= 8'h93;
  filter_in_data_log_force[3039] <= 8'h9f;
  filter_in_data_log_force[3040] <= 8'h7b;
  filter_in_data_log_force[3041] <= 8'hff;
  filter_in_data_log_force[3042] <= 8'h86;
  filter_in_data_log_force[3043] <= 8'h8e;
  filter_in_data_log_force[3044] <= 8'ha4;
  filter_in_data_log_force[3045] <= 8'h65;
  filter_in_data_log_force[3046] <= 8'hf7;
  filter_in_data_log_force[3047] <= 8'h10;
  filter_in_data_log_force[3048] <= 8'hff;
  filter_in_data_log_force[3049] <= 8'h91;
  filter_in_data_log_force[3050] <= 8'h66;
  filter_in_data_log_force[3051] <= 8'hca;
  filter_in_data_log_force[3052] <= 8'hc5;
  filter_in_data_log_force[3053] <= 8'h18;
  filter_in_data_log_force[3054] <= 8'hfa;
  filter_in_data_log_force[3055] <= 8'hde;
  filter_in_data_log_force[3056] <= 8'h28;
  filter_in_data_log_force[3057] <= 8'h70;
  filter_in_data_log_force[3058] <= 8'h1f;
  filter_in_data_log_force[3059] <= 8'hc8;
  filter_in_data_log_force[3060] <= 8'hb5;
  filter_in_data_log_force[3061] <= 8'hf0;
  filter_in_data_log_force[3062] <= 8'h87;
  filter_in_data_log_force[3063] <= 8'h60;
  filter_in_data_log_force[3064] <= 8'h1c;
  filter_in_data_log_force[3065] <= 8'hb4;
  filter_in_data_log_force[3066] <= 8'h05;
  filter_in_data_log_force[3067] <= 8'h8e;
  filter_in_data_log_force[3068] <= 8'h5d;
  filter_in_data_log_force[3069] <= 8'hf1;
  filter_in_data_log_force[3070] <= 8'h0c;
  filter_in_data_log_force[3071] <= 8'h11;
  filter_in_data_log_force[3072] <= 8'h2e;
  filter_in_data_log_force[3073] <= 8'hdf;
  filter_in_data_log_force[3074] <= 8'h94;
  filter_in_data_log_force[3075] <= 8'hf5;
  filter_in_data_log_force[3076] <= 8'h8c;
  filter_in_data_log_force[3077] <= 8'h3d;
  filter_in_data_log_force[3078] <= 8'h8a;
  filter_in_data_log_force[3079] <= 8'h74;
  filter_in_data_log_force[3080] <= 8'h3e;
  filter_in_data_log_force[3081] <= 8'h70;
  filter_in_data_log_force[3082] <= 8'h03;
  filter_in_data_log_force[3083] <= 8'hbe;
  filter_in_data_log_force[3084] <= 8'hc3;
  filter_in_data_log_force[3085] <= 8'h42;
  filter_in_data_log_force[3086] <= 8'h7e;
  filter_in_data_log_force[3087] <= 8'hdb;
  filter_in_data_log_force[3088] <= 8'h41;
  filter_in_data_log_force[3089] <= 8'h9c;
  filter_in_data_log_force[3090] <= 8'h19;
  filter_in_data_log_force[3091] <= 8'hee;
  filter_in_data_log_force[3092] <= 8'h3b;
  filter_in_data_log_force[3093] <= 8'hc3;
  filter_in_data_log_force[3094] <= 8'h98;
  filter_in_data_log_force[3095] <= 8'hf3;
  filter_in_data_log_force[3096] <= 8'h24;
  filter_in_data_log_force[3097] <= 8'ha2;
  filter_in_data_log_force[3098] <= 8'hf4;
  filter_in_data_log_force[3099] <= 8'h27;
  filter_in_data_log_force[3100] <= 8'h54;
  filter_in_data_log_force[3101] <= 8'hcf;
  filter_in_data_log_force[3102] <= 8'h00;
  filter_in_data_log_force[3103] <= 8'h00;
  filter_in_data_log_force[3104] <= 8'h00;
  filter_in_data_log_force[3105] <= 8'h00;
  filter_in_data_log_force[3106] <= 8'h00;

  // Output data for filter_out
  filter_out_expected[   0] <= 8'h03;
  filter_out_expected[   1] <= 8'h06;
  filter_out_expected[   2] <= 8'h08;
  filter_out_expected[   3] <= 8'h06;
  filter_out_expected[   4] <= 8'h03;
  filter_out_expected[   5] <= 8'h00;
  filter_out_expected[   6] <= 8'h00;
  filter_out_expected[   7] <= 8'h00;
  filter_out_expected[   8] <= 8'h00;
  filter_out_expected[   9] <= 8'h00;
  filter_out_expected[  10] <= 8'h00;
  filter_out_expected[  11] <= 8'h03;
  filter_out_expected[  12] <= 8'h09;
  filter_out_expected[  13] <= 8'h11;
  filter_out_expected[  14] <= 8'h17;
  filter_out_expected[  15] <= 8'h17;
  filter_out_expected[  16] <= 8'h11;
  filter_out_expected[  17] <= 8'h09;
  filter_out_expected[  18] <= 8'h03;
  filter_out_expected[  19] <= 8'h00;
  filter_out_expected[  20] <= 8'hfd;
  filter_out_expected[  21] <= 8'hf7;
  filter_out_expected[  22] <= 8'hef;
  filter_out_expected[  23] <= 8'he9;
  filter_out_expected[  24] <= 8'he6;
  filter_out_expected[  25] <= 8'he6;
  filter_out_expected[  26] <= 8'he6;
  filter_out_expected[  27] <= 8'he6;
  filter_out_expected[  28] <= 8'he7;
  filter_out_expected[  29] <= 8'he7;
  filter_out_expected[  30] <= 8'he7;
  filter_out_expected[  31] <= 8'he7;
  filter_out_expected[  32] <= 8'he7;
  filter_out_expected[  33] <= 8'he7;
  filter_out_expected[  34] <= 8'he7;
  filter_out_expected[  35] <= 8'he7;
  filter_out_expected[  36] <= 8'he7;
  filter_out_expected[  37] <= 8'he7;
  filter_out_expected[  38] <= 8'he7;
  filter_out_expected[  39] <= 8'he7;
  filter_out_expected[  40] <= 8'he7;
  filter_out_expected[  41] <= 8'he7;
  filter_out_expected[  42] <= 8'he7;
  filter_out_expected[  43] <= 8'he7;
  filter_out_expected[  44] <= 8'he7;
  filter_out_expected[  45] <= 8'he7;
  filter_out_expected[  46] <= 8'he7;
  filter_out_expected[  47] <= 8'he7;
  filter_out_expected[  48] <= 8'he8;
  filter_out_expected[  49] <= 8'he8;
  filter_out_expected[  50] <= 8'he8;
  filter_out_expected[  51] <= 8'he8;
  filter_out_expected[  52] <= 8'he8;
  filter_out_expected[  53] <= 8'he8;
  filter_out_expected[  54] <= 8'he8;
  filter_out_expected[  55] <= 8'he8;
  filter_out_expected[  56] <= 8'he8;
  filter_out_expected[  57] <= 8'he8;
  filter_out_expected[  58] <= 8'he8;
  filter_out_expected[  59] <= 8'he8;
  filter_out_expected[  60] <= 8'he8;
  filter_out_expected[  61] <= 8'he8;
  filter_out_expected[  62] <= 8'he8;
  filter_out_expected[  63] <= 8'he8;
  filter_out_expected[  64] <= 8'he8;
  filter_out_expected[  65] <= 8'he8;
  filter_out_expected[  66] <= 8'he8;
  filter_out_expected[  67] <= 8'he8;
  filter_out_expected[  68] <= 8'he9;
  filter_out_expected[  69] <= 8'he9;
  filter_out_expected[  70] <= 8'he9;
  filter_out_expected[  71] <= 8'he9;
  filter_out_expected[  72] <= 8'he9;
  filter_out_expected[  73] <= 8'he9;
  filter_out_expected[  74] <= 8'he9;
  filter_out_expected[  75] <= 8'he9;
  filter_out_expected[  76] <= 8'he9;
  filter_out_expected[  77] <= 8'he9;
  filter_out_expected[  78] <= 8'he9;
  filter_out_expected[  79] <= 8'he9;
  filter_out_expected[  80] <= 8'he9;
  filter_out_expected[  81] <= 8'he9;
  filter_out_expected[  82] <= 8'he9;
  filter_out_expected[  83] <= 8'he9;
  filter_out_expected[  84] <= 8'he9;
  filter_out_expected[  85] <= 8'he9;
  filter_out_expected[  86] <= 8'he9;
  filter_out_expected[  87] <= 8'he9;
  filter_out_expected[  88] <= 8'hea;
  filter_out_expected[  89] <= 8'hea;
  filter_out_expected[  90] <= 8'hea;
  filter_out_expected[  91] <= 8'hea;
  filter_out_expected[  92] <= 8'hea;
  filter_out_expected[  93] <= 8'hea;
  filter_out_expected[  94] <= 8'hea;
  filter_out_expected[  95] <= 8'hea;
  filter_out_expected[  96] <= 8'hea;
  filter_out_expected[  97] <= 8'hea;
  filter_out_expected[  98] <= 8'hea;
  filter_out_expected[  99] <= 8'hea;
  filter_out_expected[ 100] <= 8'hea;
  filter_out_expected[ 101] <= 8'hea;
  filter_out_expected[ 102] <= 8'hea;
  filter_out_expected[ 103] <= 8'hea;
  filter_out_expected[ 104] <= 8'hea;
  filter_out_expected[ 105] <= 8'hea;
  filter_out_expected[ 106] <= 8'hea;
  filter_out_expected[ 107] <= 8'hea;
  filter_out_expected[ 108] <= 8'heb;
  filter_out_expected[ 109] <= 8'heb;
  filter_out_expected[ 110] <= 8'heb;
  filter_out_expected[ 111] <= 8'heb;
  filter_out_expected[ 112] <= 8'heb;
  filter_out_expected[ 113] <= 8'heb;
  filter_out_expected[ 114] <= 8'heb;
  filter_out_expected[ 115] <= 8'heb;
  filter_out_expected[ 116] <= 8'heb;
  filter_out_expected[ 117] <= 8'heb;
  filter_out_expected[ 118] <= 8'heb;
  filter_out_expected[ 119] <= 8'heb;
  filter_out_expected[ 120] <= 8'heb;
  filter_out_expected[ 121] <= 8'heb;
  filter_out_expected[ 122] <= 8'heb;
  filter_out_expected[ 123] <= 8'heb;
  filter_out_expected[ 124] <= 8'heb;
  filter_out_expected[ 125] <= 8'heb;
  filter_out_expected[ 126] <= 8'heb;
  filter_out_expected[ 127] <= 8'heb;
  filter_out_expected[ 128] <= 8'hec;
  filter_out_expected[ 129] <= 8'hec;
  filter_out_expected[ 130] <= 8'hec;
  filter_out_expected[ 131] <= 8'hec;
  filter_out_expected[ 132] <= 8'hec;
  filter_out_expected[ 133] <= 8'hec;
  filter_out_expected[ 134] <= 8'hec;
  filter_out_expected[ 135] <= 8'hec;
  filter_out_expected[ 136] <= 8'hec;
  filter_out_expected[ 137] <= 8'hec;
  filter_out_expected[ 138] <= 8'hec;
  filter_out_expected[ 139] <= 8'hec;
  filter_out_expected[ 140] <= 8'hec;
  filter_out_expected[ 141] <= 8'hec;
  filter_out_expected[ 142] <= 8'hec;
  filter_out_expected[ 143] <= 8'hec;
  filter_out_expected[ 144] <= 8'hec;
  filter_out_expected[ 145] <= 8'hec;
  filter_out_expected[ 146] <= 8'hec;
  filter_out_expected[ 147] <= 8'hec;
  filter_out_expected[ 148] <= 8'hed;
  filter_out_expected[ 149] <= 8'hed;
  filter_out_expected[ 150] <= 8'hed;
  filter_out_expected[ 151] <= 8'hed;
  filter_out_expected[ 152] <= 8'hed;
  filter_out_expected[ 153] <= 8'hed;
  filter_out_expected[ 154] <= 8'hed;
  filter_out_expected[ 155] <= 8'hed;
  filter_out_expected[ 156] <= 8'hed;
  filter_out_expected[ 157] <= 8'hed;
  filter_out_expected[ 158] <= 8'hed;
  filter_out_expected[ 159] <= 8'hed;
  filter_out_expected[ 160] <= 8'hed;
  filter_out_expected[ 161] <= 8'hed;
  filter_out_expected[ 162] <= 8'hed;
  filter_out_expected[ 163] <= 8'hed;
  filter_out_expected[ 164] <= 8'hed;
  filter_out_expected[ 165] <= 8'hed;
  filter_out_expected[ 166] <= 8'hed;
  filter_out_expected[ 167] <= 8'hee;
  filter_out_expected[ 168] <= 8'hee;
  filter_out_expected[ 169] <= 8'hee;
  filter_out_expected[ 170] <= 8'hee;
  filter_out_expected[ 171] <= 8'hee;
  filter_out_expected[ 172] <= 8'hee;
  filter_out_expected[ 173] <= 8'hee;
  filter_out_expected[ 174] <= 8'hee;
  filter_out_expected[ 175] <= 8'hee;
  filter_out_expected[ 176] <= 8'hee;
  filter_out_expected[ 177] <= 8'hee;
  filter_out_expected[ 178] <= 8'hee;
  filter_out_expected[ 179] <= 8'hee;
  filter_out_expected[ 180] <= 8'hee;
  filter_out_expected[ 181] <= 8'hee;
  filter_out_expected[ 182] <= 8'hee;
  filter_out_expected[ 183] <= 8'hee;
  filter_out_expected[ 184] <= 8'hee;
  filter_out_expected[ 185] <= 8'hee;
  filter_out_expected[ 186] <= 8'hee;
  filter_out_expected[ 187] <= 8'hef;
  filter_out_expected[ 188] <= 8'hef;
  filter_out_expected[ 189] <= 8'hef;
  filter_out_expected[ 190] <= 8'hef;
  filter_out_expected[ 191] <= 8'hef;
  filter_out_expected[ 192] <= 8'hef;
  filter_out_expected[ 193] <= 8'hef;
  filter_out_expected[ 194] <= 8'hef;
  filter_out_expected[ 195] <= 8'hef;
  filter_out_expected[ 196] <= 8'hef;
  filter_out_expected[ 197] <= 8'hef;
  filter_out_expected[ 198] <= 8'hef;
  filter_out_expected[ 199] <= 8'hef;
  filter_out_expected[ 200] <= 8'hef;
  filter_out_expected[ 201] <= 8'hef;
  filter_out_expected[ 202] <= 8'hef;
  filter_out_expected[ 203] <= 8'hef;
  filter_out_expected[ 204] <= 8'hef;
  filter_out_expected[ 205] <= 8'hef;
  filter_out_expected[ 206] <= 8'hef;
  filter_out_expected[ 207] <= 8'hf0;
  filter_out_expected[ 208] <= 8'hf0;
  filter_out_expected[ 209] <= 8'hf0;
  filter_out_expected[ 210] <= 8'hf0;
  filter_out_expected[ 211] <= 8'hf0;
  filter_out_expected[ 212] <= 8'hf0;
  filter_out_expected[ 213] <= 8'hf0;
  filter_out_expected[ 214] <= 8'hf0;
  filter_out_expected[ 215] <= 8'hf0;
  filter_out_expected[ 216] <= 8'hf0;
  filter_out_expected[ 217] <= 8'hf0;
  filter_out_expected[ 218] <= 8'hf0;
  filter_out_expected[ 219] <= 8'hf0;
  filter_out_expected[ 220] <= 8'hf0;
  filter_out_expected[ 221] <= 8'hf0;
  filter_out_expected[ 222] <= 8'hf0;
  filter_out_expected[ 223] <= 8'hf0;
  filter_out_expected[ 224] <= 8'hf0;
  filter_out_expected[ 225] <= 8'hf0;
  filter_out_expected[ 226] <= 8'hf0;
  filter_out_expected[ 227] <= 8'hf1;
  filter_out_expected[ 228] <= 8'hf1;
  filter_out_expected[ 229] <= 8'hf1;
  filter_out_expected[ 230] <= 8'hf1;
  filter_out_expected[ 231] <= 8'hf1;
  filter_out_expected[ 232] <= 8'hf1;
  filter_out_expected[ 233] <= 8'hf1;
  filter_out_expected[ 234] <= 8'hf1;
  filter_out_expected[ 235] <= 8'hf1;
  filter_out_expected[ 236] <= 8'hf1;
  filter_out_expected[ 237] <= 8'hf1;
  filter_out_expected[ 238] <= 8'hf1;
  filter_out_expected[ 239] <= 8'hf1;
  filter_out_expected[ 240] <= 8'hf1;
  filter_out_expected[ 241] <= 8'hf1;
  filter_out_expected[ 242] <= 8'hf1;
  filter_out_expected[ 243] <= 8'hf1;
  filter_out_expected[ 244] <= 8'hf1;
  filter_out_expected[ 245] <= 8'hf1;
  filter_out_expected[ 246] <= 8'hf1;
  filter_out_expected[ 247] <= 8'hf2;
  filter_out_expected[ 248] <= 8'hf2;
  filter_out_expected[ 249] <= 8'hf2;
  filter_out_expected[ 250] <= 8'hf2;
  filter_out_expected[ 251] <= 8'hf2;
  filter_out_expected[ 252] <= 8'hf2;
  filter_out_expected[ 253] <= 8'hf2;
  filter_out_expected[ 254] <= 8'hf2;
  filter_out_expected[ 255] <= 8'hf2;
  filter_out_expected[ 256] <= 8'hf2;
  filter_out_expected[ 257] <= 8'hf2;
  filter_out_expected[ 258] <= 8'hf2;
  filter_out_expected[ 259] <= 8'hf2;
  filter_out_expected[ 260] <= 8'hf2;
  filter_out_expected[ 261] <= 8'hf2;
  filter_out_expected[ 262] <= 8'hf2;
  filter_out_expected[ 263] <= 8'hf2;
  filter_out_expected[ 264] <= 8'hf2;
  filter_out_expected[ 265] <= 8'hf2;
  filter_out_expected[ 266] <= 8'hf3;
  filter_out_expected[ 267] <= 8'hf3;
  filter_out_expected[ 268] <= 8'hf3;
  filter_out_expected[ 269] <= 8'hf3;
  filter_out_expected[ 270] <= 8'hf3;
  filter_out_expected[ 271] <= 8'hf3;
  filter_out_expected[ 272] <= 8'hf3;
  filter_out_expected[ 273] <= 8'hf3;
  filter_out_expected[ 274] <= 8'hf3;
  filter_out_expected[ 275] <= 8'hf3;
  filter_out_expected[ 276] <= 8'hf3;
  filter_out_expected[ 277] <= 8'hf3;
  filter_out_expected[ 278] <= 8'hf3;
  filter_out_expected[ 279] <= 8'hf3;
  filter_out_expected[ 280] <= 8'hf3;
  filter_out_expected[ 281] <= 8'hf3;
  filter_out_expected[ 282] <= 8'hf3;
  filter_out_expected[ 283] <= 8'hf3;
  filter_out_expected[ 284] <= 8'hf3;
  filter_out_expected[ 285] <= 8'hf3;
  filter_out_expected[ 286] <= 8'hf4;
  filter_out_expected[ 287] <= 8'hf4;
  filter_out_expected[ 288] <= 8'hf4;
  filter_out_expected[ 289] <= 8'hf4;
  filter_out_expected[ 290] <= 8'hf4;
  filter_out_expected[ 291] <= 8'hf4;
  filter_out_expected[ 292] <= 8'hf4;
  filter_out_expected[ 293] <= 8'hf4;
  filter_out_expected[ 294] <= 8'hf4;
  filter_out_expected[ 295] <= 8'hf4;
  filter_out_expected[ 296] <= 8'hf4;
  filter_out_expected[ 297] <= 8'hf4;
  filter_out_expected[ 298] <= 8'hf4;
  filter_out_expected[ 299] <= 8'hf4;
  filter_out_expected[ 300] <= 8'hf4;
  filter_out_expected[ 301] <= 8'hf4;
  filter_out_expected[ 302] <= 8'hf4;
  filter_out_expected[ 303] <= 8'hf4;
  filter_out_expected[ 304] <= 8'hf4;
  filter_out_expected[ 305] <= 8'hf4;
  filter_out_expected[ 306] <= 8'hf5;
  filter_out_expected[ 307] <= 8'hf5;
  filter_out_expected[ 308] <= 8'hf5;
  filter_out_expected[ 309] <= 8'hf5;
  filter_out_expected[ 310] <= 8'hf5;
  filter_out_expected[ 311] <= 8'hf5;
  filter_out_expected[ 312] <= 8'hf5;
  filter_out_expected[ 313] <= 8'hf5;
  filter_out_expected[ 314] <= 8'hf5;
  filter_out_expected[ 315] <= 8'hf5;
  filter_out_expected[ 316] <= 8'hf5;
  filter_out_expected[ 317] <= 8'hf5;
  filter_out_expected[ 318] <= 8'hf5;
  filter_out_expected[ 319] <= 8'hf5;
  filter_out_expected[ 320] <= 8'hf5;
  filter_out_expected[ 321] <= 8'hf5;
  filter_out_expected[ 322] <= 8'hf5;
  filter_out_expected[ 323] <= 8'hf5;
  filter_out_expected[ 324] <= 8'hf5;
  filter_out_expected[ 325] <= 8'hf5;
  filter_out_expected[ 326] <= 8'hf6;
  filter_out_expected[ 327] <= 8'hf6;
  filter_out_expected[ 328] <= 8'hf6;
  filter_out_expected[ 329] <= 8'hf6;
  filter_out_expected[ 330] <= 8'hf6;
  filter_out_expected[ 331] <= 8'hf6;
  filter_out_expected[ 332] <= 8'hf6;
  filter_out_expected[ 333] <= 8'hf6;
  filter_out_expected[ 334] <= 8'hf6;
  filter_out_expected[ 335] <= 8'hf6;
  filter_out_expected[ 336] <= 8'hf6;
  filter_out_expected[ 337] <= 8'hf6;
  filter_out_expected[ 338] <= 8'hf6;
  filter_out_expected[ 339] <= 8'hf6;
  filter_out_expected[ 340] <= 8'hf6;
  filter_out_expected[ 341] <= 8'hf6;
  filter_out_expected[ 342] <= 8'hf6;
  filter_out_expected[ 343] <= 8'hf6;
  filter_out_expected[ 344] <= 8'hf6;
  filter_out_expected[ 345] <= 8'hf6;
  filter_out_expected[ 346] <= 8'hf7;
  filter_out_expected[ 347] <= 8'hf7;
  filter_out_expected[ 348] <= 8'hf7;
  filter_out_expected[ 349] <= 8'hf7;
  filter_out_expected[ 350] <= 8'hf7;
  filter_out_expected[ 351] <= 8'hf7;
  filter_out_expected[ 352] <= 8'hf7;
  filter_out_expected[ 353] <= 8'hf7;
  filter_out_expected[ 354] <= 8'hf7;
  filter_out_expected[ 355] <= 8'hf7;
  filter_out_expected[ 356] <= 8'hf7;
  filter_out_expected[ 357] <= 8'hf7;
  filter_out_expected[ 358] <= 8'hf7;
  filter_out_expected[ 359] <= 8'hf7;
  filter_out_expected[ 360] <= 8'hf7;
  filter_out_expected[ 361] <= 8'hf7;
  filter_out_expected[ 362] <= 8'hf7;
  filter_out_expected[ 363] <= 8'hf7;
  filter_out_expected[ 364] <= 8'hf7;
  filter_out_expected[ 365] <= 8'hf8;
  filter_out_expected[ 366] <= 8'hf8;
  filter_out_expected[ 367] <= 8'hf8;
  filter_out_expected[ 368] <= 8'hf8;
  filter_out_expected[ 369] <= 8'hf8;
  filter_out_expected[ 370] <= 8'hf8;
  filter_out_expected[ 371] <= 8'hf8;
  filter_out_expected[ 372] <= 8'hf8;
  filter_out_expected[ 373] <= 8'hf8;
  filter_out_expected[ 374] <= 8'hf8;
  filter_out_expected[ 375] <= 8'hf8;
  filter_out_expected[ 376] <= 8'hf8;
  filter_out_expected[ 377] <= 8'hf8;
  filter_out_expected[ 378] <= 8'hf8;
  filter_out_expected[ 379] <= 8'hf8;
  filter_out_expected[ 380] <= 8'hf8;
  filter_out_expected[ 381] <= 8'hf8;
  filter_out_expected[ 382] <= 8'hf8;
  filter_out_expected[ 383] <= 8'hf8;
  filter_out_expected[ 384] <= 8'hf8;
  filter_out_expected[ 385] <= 8'hf9;
  filter_out_expected[ 386] <= 8'hf9;
  filter_out_expected[ 387] <= 8'hf9;
  filter_out_expected[ 388] <= 8'hf9;
  filter_out_expected[ 389] <= 8'hf9;
  filter_out_expected[ 390] <= 8'hf9;
  filter_out_expected[ 391] <= 8'hf9;
  filter_out_expected[ 392] <= 8'hf9;
  filter_out_expected[ 393] <= 8'hf9;
  filter_out_expected[ 394] <= 8'hf9;
  filter_out_expected[ 395] <= 8'hf9;
  filter_out_expected[ 396] <= 8'hf9;
  filter_out_expected[ 397] <= 8'hf9;
  filter_out_expected[ 398] <= 8'hf9;
  filter_out_expected[ 399] <= 8'hf9;
  filter_out_expected[ 400] <= 8'hf9;
  filter_out_expected[ 401] <= 8'hf9;
  filter_out_expected[ 402] <= 8'hf9;
  filter_out_expected[ 403] <= 8'hf9;
  filter_out_expected[ 404] <= 8'hf9;
  filter_out_expected[ 405] <= 8'hfa;
  filter_out_expected[ 406] <= 8'hfa;
  filter_out_expected[ 407] <= 8'hfa;
  filter_out_expected[ 408] <= 8'hfa;
  filter_out_expected[ 409] <= 8'hfa;
  filter_out_expected[ 410] <= 8'hfa;
  filter_out_expected[ 411] <= 8'hfa;
  filter_out_expected[ 412] <= 8'hfa;
  filter_out_expected[ 413] <= 8'hfa;
  filter_out_expected[ 414] <= 8'hfa;
  filter_out_expected[ 415] <= 8'hfa;
  filter_out_expected[ 416] <= 8'hfa;
  filter_out_expected[ 417] <= 8'hfa;
  filter_out_expected[ 418] <= 8'hfa;
  filter_out_expected[ 419] <= 8'hfa;
  filter_out_expected[ 420] <= 8'hfa;
  filter_out_expected[ 421] <= 8'hfa;
  filter_out_expected[ 422] <= 8'hfa;
  filter_out_expected[ 423] <= 8'hfa;
  filter_out_expected[ 424] <= 8'hfa;
  filter_out_expected[ 425] <= 8'hfb;
  filter_out_expected[ 426] <= 8'hfb;
  filter_out_expected[ 427] <= 8'hfb;
  filter_out_expected[ 428] <= 8'hfb;
  filter_out_expected[ 429] <= 8'hfb;
  filter_out_expected[ 430] <= 8'hfb;
  filter_out_expected[ 431] <= 8'hfb;
  filter_out_expected[ 432] <= 8'hfb;
  filter_out_expected[ 433] <= 8'hfb;
  filter_out_expected[ 434] <= 8'hfb;
  filter_out_expected[ 435] <= 8'hfb;
  filter_out_expected[ 436] <= 8'hfb;
  filter_out_expected[ 437] <= 8'hfb;
  filter_out_expected[ 438] <= 8'hfb;
  filter_out_expected[ 439] <= 8'hfb;
  filter_out_expected[ 440] <= 8'hfb;
  filter_out_expected[ 441] <= 8'hfb;
  filter_out_expected[ 442] <= 8'hfb;
  filter_out_expected[ 443] <= 8'hfb;
  filter_out_expected[ 444] <= 8'hfb;
  filter_out_expected[ 445] <= 8'hfc;
  filter_out_expected[ 446] <= 8'hfc;
  filter_out_expected[ 447] <= 8'hfc;
  filter_out_expected[ 448] <= 8'hfc;
  filter_out_expected[ 449] <= 8'hfc;
  filter_out_expected[ 450] <= 8'hfc;
  filter_out_expected[ 451] <= 8'hfc;
  filter_out_expected[ 452] <= 8'hfc;
  filter_out_expected[ 453] <= 8'hfc;
  filter_out_expected[ 454] <= 8'hfc;
  filter_out_expected[ 455] <= 8'hfc;
  filter_out_expected[ 456] <= 8'hfc;
  filter_out_expected[ 457] <= 8'hfc;
  filter_out_expected[ 458] <= 8'hfc;
  filter_out_expected[ 459] <= 8'hfc;
  filter_out_expected[ 460] <= 8'hfc;
  filter_out_expected[ 461] <= 8'hfc;
  filter_out_expected[ 462] <= 8'hfc;
  filter_out_expected[ 463] <= 8'hfc;
  filter_out_expected[ 464] <= 8'hfc;
  filter_out_expected[ 465] <= 8'hfd;
  filter_out_expected[ 466] <= 8'hfd;
  filter_out_expected[ 467] <= 8'hfd;
  filter_out_expected[ 468] <= 8'hfd;
  filter_out_expected[ 469] <= 8'hfd;
  filter_out_expected[ 470] <= 8'hfd;
  filter_out_expected[ 471] <= 8'hfd;
  filter_out_expected[ 472] <= 8'hfd;
  filter_out_expected[ 473] <= 8'hfd;
  filter_out_expected[ 474] <= 8'hfd;
  filter_out_expected[ 475] <= 8'hfd;
  filter_out_expected[ 476] <= 8'hfd;
  filter_out_expected[ 477] <= 8'hfd;
  filter_out_expected[ 478] <= 8'hfd;
  filter_out_expected[ 479] <= 8'hfd;
  filter_out_expected[ 480] <= 8'hfd;
  filter_out_expected[ 481] <= 8'hfd;
  filter_out_expected[ 482] <= 8'hfd;
  filter_out_expected[ 483] <= 8'hfd;
  filter_out_expected[ 484] <= 8'hfe;
  filter_out_expected[ 485] <= 8'hfe;
  filter_out_expected[ 486] <= 8'hfe;
  filter_out_expected[ 487] <= 8'hfe;
  filter_out_expected[ 488] <= 8'hfe;
  filter_out_expected[ 489] <= 8'hfe;
  filter_out_expected[ 490] <= 8'hfe;
  filter_out_expected[ 491] <= 8'hfe;
  filter_out_expected[ 492] <= 8'hfe;
  filter_out_expected[ 493] <= 8'hfe;
  filter_out_expected[ 494] <= 8'hfe;
  filter_out_expected[ 495] <= 8'hfe;
  filter_out_expected[ 496] <= 8'hfe;
  filter_out_expected[ 497] <= 8'hfe;
  filter_out_expected[ 498] <= 8'hfe;
  filter_out_expected[ 499] <= 8'hfe;
  filter_out_expected[ 500] <= 8'hfe;
  filter_out_expected[ 501] <= 8'hfe;
  filter_out_expected[ 502] <= 8'hfe;
  filter_out_expected[ 503] <= 8'hfe;
  filter_out_expected[ 504] <= 8'hff;
  filter_out_expected[ 505] <= 8'hff;
  filter_out_expected[ 506] <= 8'hff;
  filter_out_expected[ 507] <= 8'hff;
  filter_out_expected[ 508] <= 8'hff;
  filter_out_expected[ 509] <= 8'hff;
  filter_out_expected[ 510] <= 8'hff;
  filter_out_expected[ 511] <= 8'hff;
  filter_out_expected[ 512] <= 8'hff;
  filter_out_expected[ 513] <= 8'hff;
  filter_out_expected[ 514] <= 8'hff;
  filter_out_expected[ 515] <= 8'hff;
  filter_out_expected[ 516] <= 8'hff;
  filter_out_expected[ 517] <= 8'hff;
  filter_out_expected[ 518] <= 8'hff;
  filter_out_expected[ 519] <= 8'hff;
  filter_out_expected[ 520] <= 8'hff;
  filter_out_expected[ 521] <= 8'hff;
  filter_out_expected[ 522] <= 8'hff;
  filter_out_expected[ 523] <= 8'hff;
  filter_out_expected[ 524] <= 8'h00;
  filter_out_expected[ 525] <= 8'h00;
  filter_out_expected[ 526] <= 8'h00;
  filter_out_expected[ 527] <= 8'h00;
  filter_out_expected[ 528] <= 8'h00;
  filter_out_expected[ 529] <= 8'h00;
  filter_out_expected[ 530] <= 8'h00;
  filter_out_expected[ 531] <= 8'h00;
  filter_out_expected[ 532] <= 8'h00;
  filter_out_expected[ 533] <= 8'h00;
  filter_out_expected[ 534] <= 8'h00;
  filter_out_expected[ 535] <= 8'h00;
  filter_out_expected[ 536] <= 8'h00;
  filter_out_expected[ 537] <= 8'h00;
  filter_out_expected[ 538] <= 8'h00;
  filter_out_expected[ 539] <= 8'h00;
  filter_out_expected[ 540] <= 8'h00;
  filter_out_expected[ 541] <= 8'h00;
  filter_out_expected[ 542] <= 8'h00;
  filter_out_expected[ 543] <= 8'h00;
  filter_out_expected[ 544] <= 8'h01;
  filter_out_expected[ 545] <= 8'h01;
  filter_out_expected[ 546] <= 8'h01;
  filter_out_expected[ 547] <= 8'h01;
  filter_out_expected[ 548] <= 8'h01;
  filter_out_expected[ 549] <= 8'h01;
  filter_out_expected[ 550] <= 8'h01;
  filter_out_expected[ 551] <= 8'h01;
  filter_out_expected[ 552] <= 8'h01;
  filter_out_expected[ 553] <= 8'h01;
  filter_out_expected[ 554] <= 8'h01;
  filter_out_expected[ 555] <= 8'h01;
  filter_out_expected[ 556] <= 8'h01;
  filter_out_expected[ 557] <= 8'h01;
  filter_out_expected[ 558] <= 8'h01;
  filter_out_expected[ 559] <= 8'h01;
  filter_out_expected[ 560] <= 8'h01;
  filter_out_expected[ 561] <= 8'h01;
  filter_out_expected[ 562] <= 8'h01;
  filter_out_expected[ 563] <= 8'h01;
  filter_out_expected[ 564] <= 8'h02;
  filter_out_expected[ 565] <= 8'h02;
  filter_out_expected[ 566] <= 8'h02;
  filter_out_expected[ 567] <= 8'h02;
  filter_out_expected[ 568] <= 8'h02;
  filter_out_expected[ 569] <= 8'h02;
  filter_out_expected[ 570] <= 8'h02;
  filter_out_expected[ 571] <= 8'h02;
  filter_out_expected[ 572] <= 8'h02;
  filter_out_expected[ 573] <= 8'h02;
  filter_out_expected[ 574] <= 8'h02;
  filter_out_expected[ 575] <= 8'h02;
  filter_out_expected[ 576] <= 8'h02;
  filter_out_expected[ 577] <= 8'h02;
  filter_out_expected[ 578] <= 8'h02;
  filter_out_expected[ 579] <= 8'h02;
  filter_out_expected[ 580] <= 8'h02;
  filter_out_expected[ 581] <= 8'h02;
  filter_out_expected[ 582] <= 8'h02;
  filter_out_expected[ 583] <= 8'h02;
  filter_out_expected[ 584] <= 8'h03;
  filter_out_expected[ 585] <= 8'h03;
  filter_out_expected[ 586] <= 8'h03;
  filter_out_expected[ 587] <= 8'h03;
  filter_out_expected[ 588] <= 8'h03;
  filter_out_expected[ 589] <= 8'h03;
  filter_out_expected[ 590] <= 8'h03;
  filter_out_expected[ 591] <= 8'h03;
  filter_out_expected[ 592] <= 8'h03;
  filter_out_expected[ 593] <= 8'h03;
  filter_out_expected[ 594] <= 8'h03;
  filter_out_expected[ 595] <= 8'h03;
  filter_out_expected[ 596] <= 8'h03;
  filter_out_expected[ 597] <= 8'h03;
  filter_out_expected[ 598] <= 8'h03;
  filter_out_expected[ 599] <= 8'h03;
  filter_out_expected[ 600] <= 8'h03;
  filter_out_expected[ 601] <= 8'h03;
  filter_out_expected[ 602] <= 8'h03;
  filter_out_expected[ 603] <= 8'h04;
  filter_out_expected[ 604] <= 8'h04;
  filter_out_expected[ 605] <= 8'h04;
  filter_out_expected[ 606] <= 8'h04;
  filter_out_expected[ 607] <= 8'h04;
  filter_out_expected[ 608] <= 8'h04;
  filter_out_expected[ 609] <= 8'h04;
  filter_out_expected[ 610] <= 8'h04;
  filter_out_expected[ 611] <= 8'h04;
  filter_out_expected[ 612] <= 8'h04;
  filter_out_expected[ 613] <= 8'h04;
  filter_out_expected[ 614] <= 8'h04;
  filter_out_expected[ 615] <= 8'h04;
  filter_out_expected[ 616] <= 8'h04;
  filter_out_expected[ 617] <= 8'h04;
  filter_out_expected[ 618] <= 8'h04;
  filter_out_expected[ 619] <= 8'h04;
  filter_out_expected[ 620] <= 8'h04;
  filter_out_expected[ 621] <= 8'h04;
  filter_out_expected[ 622] <= 8'h04;
  filter_out_expected[ 623] <= 8'h05;
  filter_out_expected[ 624] <= 8'h05;
  filter_out_expected[ 625] <= 8'h05;
  filter_out_expected[ 626] <= 8'h05;
  filter_out_expected[ 627] <= 8'h05;
  filter_out_expected[ 628] <= 8'h05;
  filter_out_expected[ 629] <= 8'h05;
  filter_out_expected[ 630] <= 8'h05;
  filter_out_expected[ 631] <= 8'h05;
  filter_out_expected[ 632] <= 8'h05;
  filter_out_expected[ 633] <= 8'h05;
  filter_out_expected[ 634] <= 8'h05;
  filter_out_expected[ 635] <= 8'h05;
  filter_out_expected[ 636] <= 8'h05;
  filter_out_expected[ 637] <= 8'h05;
  filter_out_expected[ 638] <= 8'h05;
  filter_out_expected[ 639] <= 8'h05;
  filter_out_expected[ 640] <= 8'h05;
  filter_out_expected[ 641] <= 8'h05;
  filter_out_expected[ 642] <= 8'h05;
  filter_out_expected[ 643] <= 8'h06;
  filter_out_expected[ 644] <= 8'h06;
  filter_out_expected[ 645] <= 8'h06;
  filter_out_expected[ 646] <= 8'h06;
  filter_out_expected[ 647] <= 8'h06;
  filter_out_expected[ 648] <= 8'h06;
  filter_out_expected[ 649] <= 8'h06;
  filter_out_expected[ 650] <= 8'h06;
  filter_out_expected[ 651] <= 8'h06;
  filter_out_expected[ 652] <= 8'h06;
  filter_out_expected[ 653] <= 8'h06;
  filter_out_expected[ 654] <= 8'h06;
  filter_out_expected[ 655] <= 8'h06;
  filter_out_expected[ 656] <= 8'h06;
  filter_out_expected[ 657] <= 8'h06;
  filter_out_expected[ 658] <= 8'h06;
  filter_out_expected[ 659] <= 8'h06;
  filter_out_expected[ 660] <= 8'h06;
  filter_out_expected[ 661] <= 8'h06;
  filter_out_expected[ 662] <= 8'h06;
  filter_out_expected[ 663] <= 8'h07;
  filter_out_expected[ 664] <= 8'h07;
  filter_out_expected[ 665] <= 8'h07;
  filter_out_expected[ 666] <= 8'h07;
  filter_out_expected[ 667] <= 8'h07;
  filter_out_expected[ 668] <= 8'h07;
  filter_out_expected[ 669] <= 8'h07;
  filter_out_expected[ 670] <= 8'h07;
  filter_out_expected[ 671] <= 8'h07;
  filter_out_expected[ 672] <= 8'h07;
  filter_out_expected[ 673] <= 8'h07;
  filter_out_expected[ 674] <= 8'h07;
  filter_out_expected[ 675] <= 8'h07;
  filter_out_expected[ 676] <= 8'h07;
  filter_out_expected[ 677] <= 8'h07;
  filter_out_expected[ 678] <= 8'h07;
  filter_out_expected[ 679] <= 8'h07;
  filter_out_expected[ 680] <= 8'h07;
  filter_out_expected[ 681] <= 8'h07;
  filter_out_expected[ 682] <= 8'h07;
  filter_out_expected[ 683] <= 8'h08;
  filter_out_expected[ 684] <= 8'h08;
  filter_out_expected[ 685] <= 8'h08;
  filter_out_expected[ 686] <= 8'h08;
  filter_out_expected[ 687] <= 8'h08;
  filter_out_expected[ 688] <= 8'h08;
  filter_out_expected[ 689] <= 8'h08;
  filter_out_expected[ 690] <= 8'h08;
  filter_out_expected[ 691] <= 8'h08;
  filter_out_expected[ 692] <= 8'h08;
  filter_out_expected[ 693] <= 8'h08;
  filter_out_expected[ 694] <= 8'h08;
  filter_out_expected[ 695] <= 8'h08;
  filter_out_expected[ 696] <= 8'h08;
  filter_out_expected[ 697] <= 8'h08;
  filter_out_expected[ 698] <= 8'h08;
  filter_out_expected[ 699] <= 8'h08;
  filter_out_expected[ 700] <= 8'h08;
  filter_out_expected[ 701] <= 8'h08;
  filter_out_expected[ 702] <= 8'h08;
  filter_out_expected[ 703] <= 8'h09;
  filter_out_expected[ 704] <= 8'h09;
  filter_out_expected[ 705] <= 8'h09;
  filter_out_expected[ 706] <= 8'h09;
  filter_out_expected[ 707] <= 8'h09;
  filter_out_expected[ 708] <= 8'h09;
  filter_out_expected[ 709] <= 8'h09;
  filter_out_expected[ 710] <= 8'h09;
  filter_out_expected[ 711] <= 8'h09;
  filter_out_expected[ 712] <= 8'h09;
  filter_out_expected[ 713] <= 8'h09;
  filter_out_expected[ 714] <= 8'h09;
  filter_out_expected[ 715] <= 8'h09;
  filter_out_expected[ 716] <= 8'h09;
  filter_out_expected[ 717] <= 8'h09;
  filter_out_expected[ 718] <= 8'h09;
  filter_out_expected[ 719] <= 8'h09;
  filter_out_expected[ 720] <= 8'h09;
  filter_out_expected[ 721] <= 8'h09;
  filter_out_expected[ 722] <= 8'h0a;
  filter_out_expected[ 723] <= 8'h0a;
  filter_out_expected[ 724] <= 8'h0a;
  filter_out_expected[ 725] <= 8'h0a;
  filter_out_expected[ 726] <= 8'h0a;
  filter_out_expected[ 727] <= 8'h0a;
  filter_out_expected[ 728] <= 8'h0a;
  filter_out_expected[ 729] <= 8'h0a;
  filter_out_expected[ 730] <= 8'h0a;
  filter_out_expected[ 731] <= 8'h0a;
  filter_out_expected[ 732] <= 8'h0a;
  filter_out_expected[ 733] <= 8'h0a;
  filter_out_expected[ 734] <= 8'h0a;
  filter_out_expected[ 735] <= 8'h0a;
  filter_out_expected[ 736] <= 8'h0a;
  filter_out_expected[ 737] <= 8'h0a;
  filter_out_expected[ 738] <= 8'h0a;
  filter_out_expected[ 739] <= 8'h0a;
  filter_out_expected[ 740] <= 8'h0a;
  filter_out_expected[ 741] <= 8'h0a;
  filter_out_expected[ 742] <= 8'h0b;
  filter_out_expected[ 743] <= 8'h0b;
  filter_out_expected[ 744] <= 8'h0b;
  filter_out_expected[ 745] <= 8'h0b;
  filter_out_expected[ 746] <= 8'h0b;
  filter_out_expected[ 747] <= 8'h0b;
  filter_out_expected[ 748] <= 8'h0b;
  filter_out_expected[ 749] <= 8'h0b;
  filter_out_expected[ 750] <= 8'h0b;
  filter_out_expected[ 751] <= 8'h0b;
  filter_out_expected[ 752] <= 8'h0b;
  filter_out_expected[ 753] <= 8'h0b;
  filter_out_expected[ 754] <= 8'h0b;
  filter_out_expected[ 755] <= 8'h0b;
  filter_out_expected[ 756] <= 8'h0b;
  filter_out_expected[ 757] <= 8'h0b;
  filter_out_expected[ 758] <= 8'h0b;
  filter_out_expected[ 759] <= 8'h0b;
  filter_out_expected[ 760] <= 8'h0b;
  filter_out_expected[ 761] <= 8'h0b;
  filter_out_expected[ 762] <= 8'h0c;
  filter_out_expected[ 763] <= 8'h0c;
  filter_out_expected[ 764] <= 8'h0c;
  filter_out_expected[ 765] <= 8'h0c;
  filter_out_expected[ 766] <= 8'h0c;
  filter_out_expected[ 767] <= 8'h0c;
  filter_out_expected[ 768] <= 8'h0c;
  filter_out_expected[ 769] <= 8'h0c;
  filter_out_expected[ 770] <= 8'h0c;
  filter_out_expected[ 771] <= 8'h0c;
  filter_out_expected[ 772] <= 8'h0c;
  filter_out_expected[ 773] <= 8'h0c;
  filter_out_expected[ 774] <= 8'h0c;
  filter_out_expected[ 775] <= 8'h0c;
  filter_out_expected[ 776] <= 8'h0c;
  filter_out_expected[ 777] <= 8'h0c;
  filter_out_expected[ 778] <= 8'h0c;
  filter_out_expected[ 779] <= 8'h0c;
  filter_out_expected[ 780] <= 8'h0c;
  filter_out_expected[ 781] <= 8'h0c;
  filter_out_expected[ 782] <= 8'h0d;
  filter_out_expected[ 783] <= 8'h0d;
  filter_out_expected[ 784] <= 8'h0d;
  filter_out_expected[ 785] <= 8'h0d;
  filter_out_expected[ 786] <= 8'h0d;
  filter_out_expected[ 787] <= 8'h0d;
  filter_out_expected[ 788] <= 8'h0d;
  filter_out_expected[ 789] <= 8'h0d;
  filter_out_expected[ 790] <= 8'h0d;
  filter_out_expected[ 791] <= 8'h0d;
  filter_out_expected[ 792] <= 8'h0d;
  filter_out_expected[ 793] <= 8'h0d;
  filter_out_expected[ 794] <= 8'h0d;
  filter_out_expected[ 795] <= 8'h0d;
  filter_out_expected[ 796] <= 8'h0d;
  filter_out_expected[ 797] <= 8'h0d;
  filter_out_expected[ 798] <= 8'h0d;
  filter_out_expected[ 799] <= 8'h0d;
  filter_out_expected[ 800] <= 8'h0d;
  filter_out_expected[ 801] <= 8'h0d;
  filter_out_expected[ 802] <= 8'h0e;
  filter_out_expected[ 803] <= 8'h0e;
  filter_out_expected[ 804] <= 8'h0e;
  filter_out_expected[ 805] <= 8'h0e;
  filter_out_expected[ 806] <= 8'h0e;
  filter_out_expected[ 807] <= 8'h0e;
  filter_out_expected[ 808] <= 8'h0e;
  filter_out_expected[ 809] <= 8'h0e;
  filter_out_expected[ 810] <= 8'h0e;
  filter_out_expected[ 811] <= 8'h0e;
  filter_out_expected[ 812] <= 8'h0e;
  filter_out_expected[ 813] <= 8'h0e;
  filter_out_expected[ 814] <= 8'h0e;
  filter_out_expected[ 815] <= 8'h0e;
  filter_out_expected[ 816] <= 8'h0e;
  filter_out_expected[ 817] <= 8'h0e;
  filter_out_expected[ 818] <= 8'h0e;
  filter_out_expected[ 819] <= 8'h0e;
  filter_out_expected[ 820] <= 8'h0e;
  filter_out_expected[ 821] <= 8'h0f;
  filter_out_expected[ 822] <= 8'h0f;
  filter_out_expected[ 823] <= 8'h0f;
  filter_out_expected[ 824] <= 8'h0f;
  filter_out_expected[ 825] <= 8'h0f;
  filter_out_expected[ 826] <= 8'h0f;
  filter_out_expected[ 827] <= 8'h0f;
  filter_out_expected[ 828] <= 8'h0f;
  filter_out_expected[ 829] <= 8'h0f;
  filter_out_expected[ 830] <= 8'h0f;
  filter_out_expected[ 831] <= 8'h0f;
  filter_out_expected[ 832] <= 8'h0f;
  filter_out_expected[ 833] <= 8'h0f;
  filter_out_expected[ 834] <= 8'h0f;
  filter_out_expected[ 835] <= 8'h0f;
  filter_out_expected[ 836] <= 8'h0f;
  filter_out_expected[ 837] <= 8'h0f;
  filter_out_expected[ 838] <= 8'h0f;
  filter_out_expected[ 839] <= 8'h0f;
  filter_out_expected[ 840] <= 8'h0f;
  filter_out_expected[ 841] <= 8'h10;
  filter_out_expected[ 842] <= 8'h10;
  filter_out_expected[ 843] <= 8'h10;
  filter_out_expected[ 844] <= 8'h10;
  filter_out_expected[ 845] <= 8'h10;
  filter_out_expected[ 846] <= 8'h10;
  filter_out_expected[ 847] <= 8'h10;
  filter_out_expected[ 848] <= 8'h10;
  filter_out_expected[ 849] <= 8'h10;
  filter_out_expected[ 850] <= 8'h10;
  filter_out_expected[ 851] <= 8'h10;
  filter_out_expected[ 852] <= 8'h10;
  filter_out_expected[ 853] <= 8'h10;
  filter_out_expected[ 854] <= 8'h10;
  filter_out_expected[ 855] <= 8'h10;
  filter_out_expected[ 856] <= 8'h10;
  filter_out_expected[ 857] <= 8'h10;
  filter_out_expected[ 858] <= 8'h10;
  filter_out_expected[ 859] <= 8'h10;
  filter_out_expected[ 860] <= 8'h10;
  filter_out_expected[ 861] <= 8'h11;
  filter_out_expected[ 862] <= 8'h11;
  filter_out_expected[ 863] <= 8'h11;
  filter_out_expected[ 864] <= 8'h11;
  filter_out_expected[ 865] <= 8'h11;
  filter_out_expected[ 866] <= 8'h11;
  filter_out_expected[ 867] <= 8'h11;
  filter_out_expected[ 868] <= 8'h11;
  filter_out_expected[ 869] <= 8'h11;
  filter_out_expected[ 870] <= 8'h11;
  filter_out_expected[ 871] <= 8'h11;
  filter_out_expected[ 872] <= 8'h11;
  filter_out_expected[ 873] <= 8'h11;
  filter_out_expected[ 874] <= 8'h11;
  filter_out_expected[ 875] <= 8'h11;
  filter_out_expected[ 876] <= 8'h11;
  filter_out_expected[ 877] <= 8'h11;
  filter_out_expected[ 878] <= 8'h11;
  filter_out_expected[ 879] <= 8'h11;
  filter_out_expected[ 880] <= 8'h11;
  filter_out_expected[ 881] <= 8'h12;
  filter_out_expected[ 882] <= 8'h12;
  filter_out_expected[ 883] <= 8'h12;
  filter_out_expected[ 884] <= 8'h12;
  filter_out_expected[ 885] <= 8'h12;
  filter_out_expected[ 886] <= 8'h12;
  filter_out_expected[ 887] <= 8'h12;
  filter_out_expected[ 888] <= 8'h12;
  filter_out_expected[ 889] <= 8'h12;
  filter_out_expected[ 890] <= 8'h12;
  filter_out_expected[ 891] <= 8'h12;
  filter_out_expected[ 892] <= 8'h12;
  filter_out_expected[ 893] <= 8'h12;
  filter_out_expected[ 894] <= 8'h12;
  filter_out_expected[ 895] <= 8'h12;
  filter_out_expected[ 896] <= 8'h12;
  filter_out_expected[ 897] <= 8'h12;
  filter_out_expected[ 898] <= 8'h12;
  filter_out_expected[ 899] <= 8'h12;
  filter_out_expected[ 900] <= 8'h12;
  filter_out_expected[ 901] <= 8'h13;
  filter_out_expected[ 902] <= 8'h13;
  filter_out_expected[ 903] <= 8'h13;
  filter_out_expected[ 904] <= 8'h13;
  filter_out_expected[ 905] <= 8'h13;
  filter_out_expected[ 906] <= 8'h13;
  filter_out_expected[ 907] <= 8'h13;
  filter_out_expected[ 908] <= 8'h13;
  filter_out_expected[ 909] <= 8'h13;
  filter_out_expected[ 910] <= 8'h13;
  filter_out_expected[ 911] <= 8'h13;
  filter_out_expected[ 912] <= 8'h13;
  filter_out_expected[ 913] <= 8'h13;
  filter_out_expected[ 914] <= 8'h13;
  filter_out_expected[ 915] <= 8'h13;
  filter_out_expected[ 916] <= 8'h13;
  filter_out_expected[ 917] <= 8'h13;
  filter_out_expected[ 918] <= 8'h13;
  filter_out_expected[ 919] <= 8'h13;
  filter_out_expected[ 920] <= 8'h14;
  filter_out_expected[ 921] <= 8'h14;
  filter_out_expected[ 922] <= 8'h14;
  filter_out_expected[ 923] <= 8'h14;
  filter_out_expected[ 924] <= 8'h14;
  filter_out_expected[ 925] <= 8'h14;
  filter_out_expected[ 926] <= 8'h14;
  filter_out_expected[ 927] <= 8'h14;
  filter_out_expected[ 928] <= 8'h14;
  filter_out_expected[ 929] <= 8'h14;
  filter_out_expected[ 930] <= 8'h14;
  filter_out_expected[ 931] <= 8'h14;
  filter_out_expected[ 932] <= 8'h14;
  filter_out_expected[ 933] <= 8'h14;
  filter_out_expected[ 934] <= 8'h14;
  filter_out_expected[ 935] <= 8'h14;
  filter_out_expected[ 936] <= 8'h14;
  filter_out_expected[ 937] <= 8'h14;
  filter_out_expected[ 938] <= 8'h14;
  filter_out_expected[ 939] <= 8'h14;
  filter_out_expected[ 940] <= 8'h15;
  filter_out_expected[ 941] <= 8'h15;
  filter_out_expected[ 942] <= 8'h15;
  filter_out_expected[ 943] <= 8'h15;
  filter_out_expected[ 944] <= 8'h15;
  filter_out_expected[ 945] <= 8'h15;
  filter_out_expected[ 946] <= 8'h15;
  filter_out_expected[ 947] <= 8'h15;
  filter_out_expected[ 948] <= 8'h15;
  filter_out_expected[ 949] <= 8'h15;
  filter_out_expected[ 950] <= 8'h15;
  filter_out_expected[ 951] <= 8'h15;
  filter_out_expected[ 952] <= 8'h15;
  filter_out_expected[ 953] <= 8'h15;
  filter_out_expected[ 954] <= 8'h15;
  filter_out_expected[ 955] <= 8'h15;
  filter_out_expected[ 956] <= 8'h15;
  filter_out_expected[ 957] <= 8'h15;
  filter_out_expected[ 958] <= 8'h15;
  filter_out_expected[ 959] <= 8'h15;
  filter_out_expected[ 960] <= 8'h16;
  filter_out_expected[ 961] <= 8'h16;
  filter_out_expected[ 962] <= 8'h16;
  filter_out_expected[ 963] <= 8'h16;
  filter_out_expected[ 964] <= 8'h16;
  filter_out_expected[ 965] <= 8'h16;
  filter_out_expected[ 966] <= 8'h16;
  filter_out_expected[ 967] <= 8'h16;
  filter_out_expected[ 968] <= 8'h16;
  filter_out_expected[ 969] <= 8'h16;
  filter_out_expected[ 970] <= 8'h16;
  filter_out_expected[ 971] <= 8'h16;
  filter_out_expected[ 972] <= 8'h16;
  filter_out_expected[ 973] <= 8'h16;
  filter_out_expected[ 974] <= 8'h16;
  filter_out_expected[ 975] <= 8'h16;
  filter_out_expected[ 976] <= 8'h16;
  filter_out_expected[ 977] <= 8'h16;
  filter_out_expected[ 978] <= 8'h16;
  filter_out_expected[ 979] <= 8'h16;
  filter_out_expected[ 980] <= 8'h17;
  filter_out_expected[ 981] <= 8'h17;
  filter_out_expected[ 982] <= 8'h17;
  filter_out_expected[ 983] <= 8'h17;
  filter_out_expected[ 984] <= 8'h17;
  filter_out_expected[ 985] <= 8'h17;
  filter_out_expected[ 986] <= 8'h17;
  filter_out_expected[ 987] <= 8'h17;
  filter_out_expected[ 988] <= 8'h17;
  filter_out_expected[ 989] <= 8'h17;
  filter_out_expected[ 990] <= 8'h17;
  filter_out_expected[ 991] <= 8'h17;
  filter_out_expected[ 992] <= 8'h17;
  filter_out_expected[ 993] <= 8'h17;
  filter_out_expected[ 994] <= 8'h17;
  filter_out_expected[ 995] <= 8'h17;
  filter_out_expected[ 996] <= 8'h17;
  filter_out_expected[ 997] <= 8'h17;
  filter_out_expected[ 998] <= 8'h17;
  filter_out_expected[ 999] <= 8'h17;
  filter_out_expected[1000] <= 8'h18;
  filter_out_expected[1001] <= 8'h18;
  filter_out_expected[1002] <= 8'h18;
  filter_out_expected[1003] <= 8'h18;
  filter_out_expected[1004] <= 8'h18;
  filter_out_expected[1005] <= 8'h18;
  filter_out_expected[1006] <= 8'h18;
  filter_out_expected[1007] <= 8'h18;
  filter_out_expected[1008] <= 8'h18;
  filter_out_expected[1009] <= 8'h18;
  filter_out_expected[1010] <= 8'h18;
  filter_out_expected[1011] <= 8'h18;
  filter_out_expected[1012] <= 8'h18;
  filter_out_expected[1013] <= 8'h18;
  filter_out_expected[1014] <= 8'h18;
  filter_out_expected[1015] <= 8'h18;
  filter_out_expected[1016] <= 8'h18;
  filter_out_expected[1017] <= 8'h18;
  filter_out_expected[1018] <= 8'h18;
  filter_out_expected[1019] <= 8'h18;
  filter_out_expected[1020] <= 8'h19;
  filter_out_expected[1021] <= 8'h19;
  filter_out_expected[1022] <= 8'h19;
  filter_out_expected[1023] <= 8'h19;
  filter_out_expected[1024] <= 8'h19;
  filter_out_expected[1025] <= 8'h19;
  filter_out_expected[1026] <= 8'h19;
  filter_out_expected[1027] <= 8'h19;
  filter_out_expected[1028] <= 8'h19;
  filter_out_expected[1029] <= 8'h19;
  filter_out_expected[1030] <= 8'h19;
  filter_out_expected[1031] <= 8'h19;
  filter_out_expected[1032] <= 8'h19;
  filter_out_expected[1033] <= 8'h19;
  filter_out_expected[1034] <= 8'h19;
  filter_out_expected[1035] <= 8'h19;
  filter_out_expected[1036] <= 8'h19;
  filter_out_expected[1037] <= 8'h19;
  filter_out_expected[1038] <= 8'h19;
  filter_out_expected[1039] <= 8'h19;
  filter_out_expected[1040] <= 8'h1a;
  filter_out_expected[1041] <= 8'h1a;
  filter_out_expected[1042] <= 8'h1a;
  filter_out_expected[1043] <= 8'h1a;
  filter_out_expected[1044] <= 8'h17;
  filter_out_expected[1045] <= 8'h11;
  filter_out_expected[1046] <= 8'h09;
  filter_out_expected[1047] <= 8'h03;
  filter_out_expected[1048] <= 8'h00;
  filter_out_expected[1049] <= 8'h03;
  filter_out_expected[1050] <= 8'h09;
  filter_out_expected[1051] <= 8'h11;
  filter_out_expected[1052] <= 8'h17;
  filter_out_expected[1053] <= 8'h1a;
  filter_out_expected[1054] <= 8'h1a;
  filter_out_expected[1055] <= 8'h1a;
  filter_out_expected[1056] <= 8'h1a;
  filter_out_expected[1057] <= 8'h1a;
  filter_out_expected[1058] <= 8'h1a;
  filter_out_expected[1059] <= 8'h1a;
  filter_out_expected[1060] <= 8'h1a;
  filter_out_expected[1061] <= 8'h1a;
  filter_out_expected[1062] <= 8'h19;
  filter_out_expected[1063] <= 8'h19;
  filter_out_expected[1064] <= 8'h19;
  filter_out_expected[1065] <= 8'h19;
  filter_out_expected[1066] <= 8'h18;
  filter_out_expected[1067] <= 8'h18;
  filter_out_expected[1068] <= 8'h17;
  filter_out_expected[1069] <= 8'h17;
  filter_out_expected[1070] <= 8'h16;
  filter_out_expected[1071] <= 8'h15;
  filter_out_expected[1072] <= 8'h14;
  filter_out_expected[1073] <= 8'h13;
  filter_out_expected[1074] <= 8'h12;
  filter_out_expected[1075] <= 8'h11;
  filter_out_expected[1076] <= 8'h0f;
  filter_out_expected[1077] <= 8'h0d;
  filter_out_expected[1078] <= 8'h0c;
  filter_out_expected[1079] <= 8'h0a;
  filter_out_expected[1080] <= 8'h08;
  filter_out_expected[1081] <= 8'h05;
  filter_out_expected[1082] <= 8'h03;
  filter_out_expected[1083] <= 8'h01;
  filter_out_expected[1084] <= 8'hfe;
  filter_out_expected[1085] <= 8'hfc;
  filter_out_expected[1086] <= 8'hf9;
  filter_out_expected[1087] <= 8'hf7;
  filter_out_expected[1088] <= 8'hf4;
  filter_out_expected[1089] <= 8'hf2;
  filter_out_expected[1090] <= 8'hef;
  filter_out_expected[1091] <= 8'hed;
  filter_out_expected[1092] <= 8'heb;
  filter_out_expected[1093] <= 8'he9;
  filter_out_expected[1094] <= 8'he8;
  filter_out_expected[1095] <= 8'he7;
  filter_out_expected[1096] <= 8'he7;
  filter_out_expected[1097] <= 8'he7;
  filter_out_expected[1098] <= 8'he7;
  filter_out_expected[1099] <= 8'he8;
  filter_out_expected[1100] <= 8'he9;
  filter_out_expected[1101] <= 8'heb;
  filter_out_expected[1102] <= 8'hee;
  filter_out_expected[1103] <= 8'hf1;
  filter_out_expected[1104] <= 8'hf4;
  filter_out_expected[1105] <= 8'hf8;
  filter_out_expected[1106] <= 8'hfc;
  filter_out_expected[1107] <= 8'h00;
  filter_out_expected[1108] <= 8'h04;
  filter_out_expected[1109] <= 8'h09;
  filter_out_expected[1110] <= 8'h0d;
  filter_out_expected[1111] <= 8'h10;
  filter_out_expected[1112] <= 8'h14;
  filter_out_expected[1113] <= 8'h16;
  filter_out_expected[1114] <= 8'h18;
  filter_out_expected[1115] <= 8'h19;
  filter_out_expected[1116] <= 8'h19;
  filter_out_expected[1117] <= 8'h18;
  filter_out_expected[1118] <= 8'h16;
  filter_out_expected[1119] <= 8'h14;
  filter_out_expected[1120] <= 8'h10;
  filter_out_expected[1121] <= 8'h0c;
  filter_out_expected[1122] <= 8'h07;
  filter_out_expected[1123] <= 8'h01;
  filter_out_expected[1124] <= 8'hfc;
  filter_out_expected[1125] <= 8'hf7;
  filter_out_expected[1126] <= 8'hf2;
  filter_out_expected[1127] <= 8'hee;
  filter_out_expected[1128] <= 8'hea;
  filter_out_expected[1129] <= 8'he8;
  filter_out_expected[1130] <= 8'he7;
  filter_out_expected[1131] <= 8'he8;
  filter_out_expected[1132] <= 8'hea;
  filter_out_expected[1133] <= 8'hed;
  filter_out_expected[1134] <= 8'hf2;
  filter_out_expected[1135] <= 8'hf7;
  filter_out_expected[1136] <= 8'hfd;
  filter_out_expected[1137] <= 8'h03;
  filter_out_expected[1138] <= 8'h09;
  filter_out_expected[1139] <= 8'h0f;
  filter_out_expected[1140] <= 8'h14;
  filter_out_expected[1141] <= 8'h17;
  filter_out_expected[1142] <= 8'h18;
  filter_out_expected[1143] <= 8'h18;
  filter_out_expected[1144] <= 8'h16;
  filter_out_expected[1145] <= 8'h12;
  filter_out_expected[1146] <= 8'h0d;
  filter_out_expected[1147] <= 8'h06;
  filter_out_expected[1148] <= 8'hff;
  filter_out_expected[1149] <= 8'hf8;
  filter_out_expected[1150] <= 8'hf2;
  filter_out_expected[1151] <= 8'hed;
  filter_out_expected[1152] <= 8'he9;
  filter_out_expected[1153] <= 8'he8;
  filter_out_expected[1154] <= 8'he9;
  filter_out_expected[1155] <= 8'hec;
  filter_out_expected[1156] <= 8'hf1;
  filter_out_expected[1157] <= 8'hf7;
  filter_out_expected[1158] <= 8'hff;
  filter_out_expected[1159] <= 8'h07;
  filter_out_expected[1160] <= 8'h0e;
  filter_out_expected[1161] <= 8'h13;
  filter_out_expected[1162] <= 8'h17;
  filter_out_expected[1163] <= 8'h18;
  filter_out_expected[1164] <= 8'h16;
  filter_out_expected[1165] <= 8'h12;
  filter_out_expected[1166] <= 8'h0c;
  filter_out_expected[1167] <= 8'h04;
  filter_out_expected[1168] <= 8'hfc;
  filter_out_expected[1169] <= 8'hf4;
  filter_out_expected[1170] <= 8'hee;
  filter_out_expected[1171] <= 8'hea;
  filter_out_expected[1172] <= 8'he9;
  filter_out_expected[1173] <= 8'hea;
  filter_out_expected[1174] <= 8'hef;
  filter_out_expected[1175] <= 8'hf6;
  filter_out_expected[1176] <= 8'hff;
  filter_out_expected[1177] <= 8'h08;
  filter_out_expected[1178] <= 8'h0f;
  filter_out_expected[1179] <= 8'h15;
  filter_out_expected[1180] <= 8'h17;
  filter_out_expected[1181] <= 8'h16;
  filter_out_expected[1182] <= 8'h12;
  filter_out_expected[1183] <= 8'h0b;
  filter_out_expected[1184] <= 8'h02;
  filter_out_expected[1185] <= 8'hf9;
  filter_out_expected[1186] <= 8'hf1;
  filter_out_expected[1187] <= 8'heb;
  filter_out_expected[1188] <= 8'he9;
  filter_out_expected[1189] <= 8'heb;
  filter_out_expected[1190] <= 8'hf0;
  filter_out_expected[1191] <= 8'hf8;
  filter_out_expected[1192] <= 8'h02;
  filter_out_expected[1193] <= 8'h0b;
  filter_out_expected[1194] <= 8'h12;
  filter_out_expected[1195] <= 8'h16;
  filter_out_expected[1196] <= 8'h16;
  filter_out_expected[1197] <= 8'h12;
  filter_out_expected[1198] <= 8'h0a;
  filter_out_expected[1199] <= 8'h01;
  filter_out_expected[1200] <= 8'hf7;
  filter_out_expected[1201] <= 8'hef;
  filter_out_expected[1202] <= 8'hea;
  filter_out_expected[1203] <= 8'hea;
  filter_out_expected[1204] <= 8'hef;
  filter_out_expected[1205] <= 8'hf7;
  filter_out_expected[1206] <= 8'h01;
  filter_out_expected[1207] <= 8'h0a;
  filter_out_expected[1208] <= 8'h12;
  filter_out_expected[1209] <= 8'h16;
  filter_out_expected[1210] <= 8'h15;
  filter_out_expected[1211] <= 8'h0f;
  filter_out_expected[1212] <= 8'h06;
  filter_out_expected[1213] <= 8'hfb;
  filter_out_expected[1214] <= 8'hf2;
  filter_out_expected[1215] <= 8'hec;
  filter_out_expected[1216] <= 8'heb;
  filter_out_expected[1217] <= 8'hef;
  filter_out_expected[1218] <= 8'hf7;
  filter_out_expected[1219] <= 8'h01;
  filter_out_expected[1220] <= 8'h0c;
  filter_out_expected[1221] <= 8'h13;
  filter_out_expected[1222] <= 8'h15;
  filter_out_expected[1223] <= 8'h12;
  filter_out_expected[1224] <= 8'h0a;
  filter_out_expected[1225] <= 8'h00;
  filter_out_expected[1226] <= 8'hf5;
  filter_out_expected[1227] <= 8'hee;
  filter_out_expected[1228] <= 8'heb;
  filter_out_expected[1229] <= 8'hee;
  filter_out_expected[1230] <= 8'hf6;
  filter_out_expected[1231] <= 8'h01;
  filter_out_expected[1232] <= 8'h0c;
  filter_out_expected[1233] <= 8'h13;
  filter_out_expected[1234] <= 8'h15;
  filter_out_expected[1235] <= 8'h10;
  filter_out_expected[1236] <= 8'h07;
  filter_out_expected[1237] <= 8'hfb;
  filter_out_expected[1238] <= 8'hf2;
  filter_out_expected[1239] <= 8'hec;
  filter_out_expected[1240] <= 8'hed;
  filter_out_expected[1241] <= 8'hf4;
  filter_out_expected[1242] <= 8'hfe;
  filter_out_expected[1243] <= 8'h0a;
  filter_out_expected[1244] <= 8'h12;
  filter_out_expected[1245] <= 8'h14;
  filter_out_expected[1246] <= 8'h10;
  filter_out_expected[1247] <= 8'h06;
  filter_out_expected[1248] <= 8'hfa;
  filter_out_expected[1249] <= 8'hf1;
  filter_out_expected[1250] <= 8'hec;
  filter_out_expected[1251] <= 8'hef;
  filter_out_expected[1252] <= 8'hf7;
  filter_out_expected[1253] <= 8'h03;
  filter_out_expected[1254] <= 8'h0d;
  filter_out_expected[1255] <= 8'h13;
  filter_out_expected[1256] <= 8'h12;
  filter_out_expected[1257] <= 8'h0a;
  filter_out_expected[1258] <= 8'hff;
  filter_out_expected[1259] <= 8'hf4;
  filter_out_expected[1260] <= 8'hed;
  filter_out_expected[1261] <= 8'hee;
  filter_out_expected[1262] <= 8'hf6;
  filter_out_expected[1263] <= 8'h02;
  filter_out_expected[1264] <= 8'h0d;
  filter_out_expected[1265] <= 8'h13;
  filter_out_expected[1266] <= 8'h11;
  filter_out_expected[1267] <= 8'h09;
  filter_out_expected[1268] <= 8'hfd;
  filter_out_expected[1269] <= 8'hf2;
  filter_out_expected[1270] <= 8'hed;
  filter_out_expected[1271] <= 8'hf0;
  filter_out_expected[1272] <= 8'hfa;
  filter_out_expected[1273] <= 8'h06;
  filter_out_expected[1274] <= 8'h10;
  filter_out_expected[1275] <= 8'h12;
  filter_out_expected[1276] <= 8'h0d;
  filter_out_expected[1277] <= 8'h02;
  filter_out_expected[1278] <= 8'hf6;
  filter_out_expected[1279] <= 8'hef;
  filter_out_expected[1280] <= 8'hef;
  filter_out_expected[1281] <= 8'hf7;
  filter_out_expected[1282] <= 8'h03;
  filter_out_expected[1283] <= 8'h0e;
  filter_out_expected[1284] <= 8'h12;
  filter_out_expected[1285] <= 8'h0d;
  filter_out_expected[1286] <= 8'h03;
  filter_out_expected[1287] <= 8'hf7;
  filter_out_expected[1288] <= 8'hef;
  filter_out_expected[1289] <= 8'hf0;
  filter_out_expected[1290] <= 8'hf9;
  filter_out_expected[1291] <= 8'h05;
  filter_out_expected[1292] <= 8'h0f;
  filter_out_expected[1293] <= 8'h11;
  filter_out_expected[1294] <= 8'h0b;
  filter_out_expected[1295] <= 8'hff;
  filter_out_expected[1296] <= 8'hf4;
  filter_out_expected[1297] <= 8'hef;
  filter_out_expected[1298] <= 8'hf3;
  filter_out_expected[1299] <= 8'hfe;
  filter_out_expected[1300] <= 8'h0a;
  filter_out_expected[1301] <= 8'h11;
  filter_out_expected[1302] <= 8'h0e;
  filter_out_expected[1303] <= 8'h04;
  filter_out_expected[1304] <= 8'hf8;
  filter_out_expected[1305] <= 8'hf0;
  filter_out_expected[1306] <= 8'hf1;
  filter_out_expected[1307] <= 8'hfa;
  filter_out_expected[1308] <= 8'h07;
  filter_out_expected[1309] <= 8'h0f;
  filter_out_expected[1310] <= 8'h0f;
  filter_out_expected[1311] <= 8'h06;
  filter_out_expected[1312] <= 8'hfa;
  filter_out_expected[1313] <= 8'hf1;
  filter_out_expected[1314] <= 8'hf1;
  filter_out_expected[1315] <= 8'hfa;
  filter_out_expected[1316] <= 8'h07;
  filter_out_expected[1317] <= 8'h0f;
  filter_out_expected[1318] <= 8'h0e;
  filter_out_expected[1319] <= 8'h05;
  filter_out_expected[1320] <= 8'hf8;
  filter_out_expected[1321] <= 8'hf1;
  filter_out_expected[1322] <= 8'hf3;
  filter_out_expected[1323] <= 8'hfd;
  filter_out_expected[1324] <= 8'h09;
  filter_out_expected[1325] <= 8'h0f;
  filter_out_expected[1326] <= 8'h0c;
  filter_out_expected[1327] <= 8'h01;
  filter_out_expected[1328] <= 8'hf5;
  filter_out_expected[1329] <= 8'hf1;
  filter_out_expected[1330] <= 8'hf7;
  filter_out_expected[1331] <= 8'h02;
  filter_out_expected[1332] <= 8'h0d;
  filter_out_expected[1333] <= 8'h0e;
  filter_out_expected[1334] <= 8'h06;
  filter_out_expected[1335] <= 8'hfa;
  filter_out_expected[1336] <= 8'hf2;
  filter_out_expected[1337] <= 8'hf4;
  filter_out_expected[1338] <= 8'hfe;
  filter_out_expected[1339] <= 8'h09;
  filter_out_expected[1340] <= 8'h0e;
  filter_out_expected[1341] <= 8'h09;
  filter_out_expected[1342] <= 8'hfd;
  filter_out_expected[1343] <= 8'hf4;
  filter_out_expected[1344] <= 8'hf3;
  filter_out_expected[1345] <= 8'hfc;
  filter_out_expected[1346] <= 8'h08;
  filter_out_expected[1347] <= 8'h0e;
  filter_out_expected[1348] <= 8'h0a;
  filter_out_expected[1349] <= 8'hfe;
  filter_out_expected[1350] <= 8'hf4;
  filter_out_expected[1351] <= 8'hf3;
  filter_out_expected[1352] <= 8'hfc;
  filter_out_expected[1353] <= 8'h07;
  filter_out_expected[1354] <= 8'h0d;
  filter_out_expected[1355] <= 8'h09;
  filter_out_expected[1356] <= 8'hfe;
  filter_out_expected[1357] <= 8'hf4;
  filter_out_expected[1358] <= 8'hf4;
  filter_out_expected[1359] <= 8'hfd;
  filter_out_expected[1360] <= 8'h09;
  filter_out_expected[1361] <= 8'h0d;
  filter_out_expected[1362] <= 8'h07;
  filter_out_expected[1363] <= 8'hfb;
  filter_out_expected[1364] <= 8'hf3;
  filter_out_expected[1365] <= 8'hf6;
  filter_out_expected[1366] <= 8'h01;
  filter_out_expected[1367] <= 8'h0b;
  filter_out_expected[1368] <= 8'h0c;
  filter_out_expected[1369] <= 8'h02;
  filter_out_expected[1370] <= 8'hf7;
  filter_out_expected[1371] <= 8'hf4;
  filter_out_expected[1372] <= 8'hfb;
  filter_out_expected[1373] <= 8'h06;
  filter_out_expected[1374] <= 8'h0c;
  filter_out_expected[1375] <= 8'h08;
  filter_out_expected[1376] <= 8'hfd;
  filter_out_expected[1377] <= 8'hf5;
  filter_out_expected[1378] <= 8'hf7;
  filter_out_expected[1379] <= 8'h01;
  filter_out_expected[1380] <= 8'h0a;
  filter_out_expected[1381] <= 8'h0a;
  filter_out_expected[1382] <= 8'h01;
  filter_out_expected[1383] <= 8'hf7;
  filter_out_expected[1384] <= 8'hf5;
  filter_out_expected[1385] <= 8'hfe;
  filter_out_expected[1386] <= 8'h08;
  filter_out_expected[1387] <= 8'h0b;
  filter_out_expected[1388] <= 8'h04;
  filter_out_expected[1389] <= 8'hf9;
  filter_out_expected[1390] <= 8'hf5;
  filter_out_expected[1391] <= 8'hfc;
  filter_out_expected[1392] <= 8'h06;
  filter_out_expected[1393] <= 8'h0b;
  filter_out_expected[1394] <= 8'h05;
  filter_out_expected[1395] <= 8'hfa;
  filter_out_expected[1396] <= 8'hf5;
  filter_out_expected[1397] <= 8'hfb;
  filter_out_expected[1398] <= 8'h06;
  filter_out_expected[1399] <= 8'h0b;
  filter_out_expected[1400] <= 8'h05;
  filter_out_expected[1401] <= 8'hfa;
  filter_out_expected[1402] <= 8'hf6;
  filter_out_expected[1403] <= 8'hfb;
  filter_out_expected[1404] <= 8'h06;
  filter_out_expected[1405] <= 8'h0a;
  filter_out_expected[1406] <= 8'h04;
  filter_out_expected[1407] <= 8'hfa;
  filter_out_expected[1408] <= 8'hf6;
  filter_out_expected[1409] <= 8'hfd;
  filter_out_expected[1410] <= 8'h07;
  filter_out_expected[1411] <= 8'h0a;
  filter_out_expected[1412] <= 8'h02;
  filter_out_expected[1413] <= 8'hf9;
  filter_out_expected[1414] <= 8'hf7;
  filter_out_expected[1415] <= 8'hff;
  filter_out_expected[1416] <= 8'h08;
  filter_out_expected[1417] <= 8'h08;
  filter_out_expected[1418] <= 8'h00;
  filter_out_expected[1419] <= 8'hf7;
  filter_out_expected[1420] <= 8'hf9;
  filter_out_expected[1421] <= 8'h02;
  filter_out_expected[1422] <= 8'h09;
  filter_out_expected[1423] <= 8'h06;
  filter_out_expected[1424] <= 8'hfc;
  filter_out_expected[1425] <= 8'hf7;
  filter_out_expected[1426] <= 8'hfc;
  filter_out_expected[1427] <= 8'h06;
  filter_out_expected[1428] <= 8'h09;
  filter_out_expected[1429] <= 8'h02;
  filter_out_expected[1430] <= 8'hf9;
  filter_out_expected[1431] <= 8'hf8;
  filter_out_expected[1432] <= 8'h01;
  filter_out_expected[1433] <= 8'h08;
  filter_out_expected[1434] <= 8'h06;
  filter_out_expected[1435] <= 8'hfd;
  filter_out_expected[1436] <= 8'hf8;
  filter_out_expected[1437] <= 8'hfd;
  filter_out_expected[1438] <= 8'h06;
  filter_out_expected[1439] <= 8'h08;
  filter_out_expected[1440] <= 8'h01;
  filter_out_expected[1441] <= 8'hf9;
  filter_out_expected[1442] <= 8'hfa;
  filter_out_expected[1443] <= 8'h02;
  filter_out_expected[1444] <= 8'h08;
  filter_out_expected[1445] <= 8'h03;
  filter_out_expected[1446] <= 8'hfb;
  filter_out_expected[1447] <= 8'hf9;
  filter_out_expected[1448] <= 8'h00;
  filter_out_expected[1449] <= 8'h07;
  filter_out_expected[1450] <= 8'h05;
  filter_out_expected[1451] <= 8'hfd;
  filter_out_expected[1452] <= 8'hf9;
  filter_out_expected[1453] <= 8'hfe;
  filter_out_expected[1454] <= 8'h06;
  filter_out_expected[1455] <= 8'h06;
  filter_out_expected[1456] <= 8'hff;
  filter_out_expected[1457] <= 8'hf9;
  filter_out_expected[1458] <= 8'hfd;
  filter_out_expected[1459] <= 8'h05;
  filter_out_expected[1460] <= 8'h06;
  filter_out_expected[1461] <= 8'h00;
  filter_out_expected[1462] <= 8'hf9;
  filter_out_expected[1463] <= 8'hfc;
  filter_out_expected[1464] <= 8'h04;
  filter_out_expected[1465] <= 8'h06;
  filter_out_expected[1466] <= 8'h00;
  filter_out_expected[1467] <= 8'hfa;
  filter_out_expected[1468] <= 8'hfc;
  filter_out_expected[1469] <= 8'h04;
  filter_out_expected[1470] <= 8'h06;
  filter_out_expected[1471] <= 8'h00;
  filter_out_expected[1472] <= 8'hfa;
  filter_out_expected[1473] <= 8'hfc;
  filter_out_expected[1474] <= 8'h04;
  filter_out_expected[1475] <= 8'h06;
  filter_out_expected[1476] <= 8'h00;
  filter_out_expected[1477] <= 8'hfa;
  filter_out_expected[1478] <= 8'hfd;
  filter_out_expected[1479] <= 8'h04;
  filter_out_expected[1480] <= 8'h05;
  filter_out_expected[1481] <= 8'hff;
  filter_out_expected[1482] <= 8'hfa;
  filter_out_expected[1483] <= 8'hfe;
  filter_out_expected[1484] <= 8'h05;
  filter_out_expected[1485] <= 8'h04;
  filter_out_expected[1486] <= 8'hfe;
  filter_out_expected[1487] <= 8'hfb;
  filter_out_expected[1488] <= 8'hff;
  filter_out_expected[1489] <= 8'h05;
  filter_out_expected[1490] <= 8'h03;
  filter_out_expected[1491] <= 8'hfd;
  filter_out_expected[1492] <= 8'hfb;
  filter_out_expected[1493] <= 8'h01;
  filter_out_expected[1494] <= 8'h05;
  filter_out_expected[1495] <= 8'h01;
  filter_out_expected[1496] <= 8'hfc;
  filter_out_expected[1497] <= 8'hfd;
  filter_out_expected[1498] <= 8'h03;
  filter_out_expected[1499] <= 8'h04;
  filter_out_expected[1500] <= 8'hff;
  filter_out_expected[1501] <= 8'hfb;
  filter_out_expected[1502] <= 8'hff;
  filter_out_expected[1503] <= 8'h04;
  filter_out_expected[1504] <= 8'h03;
  filter_out_expected[1505] <= 8'hfd;
  filter_out_expected[1506] <= 8'hfc;
  filter_out_expected[1507] <= 8'h01;
  filter_out_expected[1508] <= 8'h04;
  filter_out_expected[1509] <= 8'h00;
  filter_out_expected[1510] <= 8'hfc;
  filter_out_expected[1511] <= 8'hfe;
  filter_out_expected[1512] <= 8'h03;
  filter_out_expected[1513] <= 8'h03;
  filter_out_expected[1514] <= 8'hfe;
  filter_out_expected[1515] <= 8'hfc;
  filter_out_expected[1516] <= 8'h01;
  filter_out_expected[1517] <= 8'h04;
  filter_out_expected[1518] <= 8'h00;
  filter_out_expected[1519] <= 8'hfc;
  filter_out_expected[1520] <= 8'hfe;
  filter_out_expected[1521] <= 8'h03;
  filter_out_expected[1522] <= 8'h03;
  filter_out_expected[1523] <= 8'hfe;
  filter_out_expected[1524] <= 8'hfd;
  filter_out_expected[1525] <= 8'h01;
  filter_out_expected[1526] <= 8'h03;
  filter_out_expected[1527] <= 8'h00;
  filter_out_expected[1528] <= 8'hfd;
  filter_out_expected[1529] <= 8'hff;
  filter_out_expected[1530] <= 8'h03;
  filter_out_expected[1531] <= 8'h01;
  filter_out_expected[1532] <= 8'hfd;
  filter_out_expected[1533] <= 8'hfe;
  filter_out_expected[1534] <= 8'h02;
  filter_out_expected[1535] <= 8'h02;
  filter_out_expected[1536] <= 8'hfe;
  filter_out_expected[1537] <= 8'hfd;
  filter_out_expected[1538] <= 8'h01;
  filter_out_expected[1539] <= 8'h03;
  filter_out_expected[1540] <= 8'h00;
  filter_out_expected[1541] <= 8'hfd;
  filter_out_expected[1542] <= 8'h00;
  filter_out_expected[1543] <= 8'h03;
  filter_out_expected[1544] <= 8'h01;
  filter_out_expected[1545] <= 8'hfe;
  filter_out_expected[1546] <= 8'hff;
  filter_out_expected[1547] <= 8'h02;
  filter_out_expected[1548] <= 8'h01;
  filter_out_expected[1549] <= 8'hfe;
  filter_out_expected[1550] <= 8'hfe;
  filter_out_expected[1551] <= 8'h02;
  filter_out_expected[1552] <= 8'h02;
  filter_out_expected[1553] <= 8'hff;
  filter_out_expected[1554] <= 8'hfe;
  filter_out_expected[1555] <= 8'h01;
  filter_out_expected[1556] <= 8'h02;
  filter_out_expected[1557] <= 8'hff;
  filter_out_expected[1558] <= 8'hfe;
  filter_out_expected[1559] <= 8'h01;
  filter_out_expected[1560] <= 8'h02;
  filter_out_expected[1561] <= 8'h00;
  filter_out_expected[1562] <= 8'hfe;
  filter_out_expected[1563] <= 8'h00;
  filter_out_expected[1564] <= 8'h02;
  filter_out_expected[1565] <= 8'h00;
  filter_out_expected[1566] <= 8'hfe;
  filter_out_expected[1567] <= 8'h00;
  filter_out_expected[1568] <= 8'h02;
  filter_out_expected[1569] <= 8'h00;
  filter_out_expected[1570] <= 8'hfe;
  filter_out_expected[1571] <= 8'h00;
  filter_out_expected[1572] <= 8'h02;
  filter_out_expected[1573] <= 8'h00;
  filter_out_expected[1574] <= 8'hfe;
  filter_out_expected[1575] <= 8'h00;
  filter_out_expected[1576] <= 8'h01;
  filter_out_expected[1577] <= 8'h00;
  filter_out_expected[1578] <= 8'hff;
  filter_out_expected[1579] <= 8'h00;
  filter_out_expected[1580] <= 8'h01;
  filter_out_expected[1581] <= 8'h00;
  filter_out_expected[1582] <= 8'hff;
  filter_out_expected[1583] <= 8'h00;
  filter_out_expected[1584] <= 8'h01;
  filter_out_expected[1585] <= 8'h00;
  filter_out_expected[1586] <= 8'hff;
  filter_out_expected[1587] <= 8'h00;
  filter_out_expected[1588] <= 8'h01;
  filter_out_expected[1589] <= 8'h00;
  filter_out_expected[1590] <= 8'hff;
  filter_out_expected[1591] <= 8'h00;
  filter_out_expected[1592] <= 8'h01;
  filter_out_expected[1593] <= 8'h00;
  filter_out_expected[1594] <= 8'hff;
  filter_out_expected[1595] <= 8'h00;
  filter_out_expected[1596] <= 8'h01;
  filter_out_expected[1597] <= 8'hff;
  filter_out_expected[1598] <= 8'h00;
  filter_out_expected[1599] <= 8'h00;
  filter_out_expected[1600] <= 8'h00;
  filter_out_expected[1601] <= 8'hff;
  filter_out_expected[1602] <= 8'h00;
  filter_out_expected[1603] <= 8'h00;
  filter_out_expected[1604] <= 8'h00;
  filter_out_expected[1605] <= 8'h00;
  filter_out_expected[1606] <= 8'h00;
  filter_out_expected[1607] <= 8'h00;
  filter_out_expected[1608] <= 8'h00;
  filter_out_expected[1609] <= 8'h00;
  filter_out_expected[1610] <= 8'h00;
  filter_out_expected[1611] <= 8'h00;
  filter_out_expected[1612] <= 8'h00;
  filter_out_expected[1613] <= 8'h00;
  filter_out_expected[1614] <= 8'h00;
  filter_out_expected[1615] <= 8'h00;
  filter_out_expected[1616] <= 8'h00;
  filter_out_expected[1617] <= 8'h00;
  filter_out_expected[1618] <= 8'h00;
  filter_out_expected[1619] <= 8'h00;
  filter_out_expected[1620] <= 8'h00;
  filter_out_expected[1621] <= 8'h00;
  filter_out_expected[1622] <= 8'h00;
  filter_out_expected[1623] <= 8'h00;
  filter_out_expected[1624] <= 8'h00;
  filter_out_expected[1625] <= 8'h00;
  filter_out_expected[1626] <= 8'h00;
  filter_out_expected[1627] <= 8'h00;
  filter_out_expected[1628] <= 8'h00;
  filter_out_expected[1629] <= 8'h00;
  filter_out_expected[1630] <= 8'h00;
  filter_out_expected[1631] <= 8'h00;
  filter_out_expected[1632] <= 8'h00;
  filter_out_expected[1633] <= 8'h00;
  filter_out_expected[1634] <= 8'h00;
  filter_out_expected[1635] <= 8'h00;
  filter_out_expected[1636] <= 8'h00;
  filter_out_expected[1637] <= 8'h00;
  filter_out_expected[1638] <= 8'h00;
  filter_out_expected[1639] <= 8'h00;
  filter_out_expected[1640] <= 8'h00;
  filter_out_expected[1641] <= 8'h00;
  filter_out_expected[1642] <= 8'h00;
  filter_out_expected[1643] <= 8'h00;
  filter_out_expected[1644] <= 8'h00;
  filter_out_expected[1645] <= 8'h01;
  filter_out_expected[1646] <= 8'h00;
  filter_out_expected[1647] <= 8'hff;
  filter_out_expected[1648] <= 8'h00;
  filter_out_expected[1649] <= 8'h00;
  filter_out_expected[1650] <= 8'hff;
  filter_out_expected[1651] <= 8'h00;
  filter_out_expected[1652] <= 8'h01;
  filter_out_expected[1653] <= 8'h00;
  filter_out_expected[1654] <= 8'hff;
  filter_out_expected[1655] <= 8'h01;
  filter_out_expected[1656] <= 8'h00;
  filter_out_expected[1657] <= 8'hff;
  filter_out_expected[1658] <= 8'h00;
  filter_out_expected[1659] <= 8'h01;
  filter_out_expected[1660] <= 8'h00;
  filter_out_expected[1661] <= 8'hff;
  filter_out_expected[1662] <= 8'h01;
  filter_out_expected[1663] <= 8'h00;
  filter_out_expected[1664] <= 8'hff;
  filter_out_expected[1665] <= 8'h00;
  filter_out_expected[1666] <= 8'h01;
  filter_out_expected[1667] <= 8'hff;
  filter_out_expected[1668] <= 8'h00;
  filter_out_expected[1669] <= 8'h01;
  filter_out_expected[1670] <= 8'h00;
  filter_out_expected[1671] <= 8'hff;
  filter_out_expected[1672] <= 8'h01;
  filter_out_expected[1673] <= 8'h01;
  filter_out_expected[1674] <= 8'hff;
  filter_out_expected[1675] <= 8'h00;
  filter_out_expected[1676] <= 8'h01;
  filter_out_expected[1677] <= 8'hff;
  filter_out_expected[1678] <= 8'hff;
  filter_out_expected[1679] <= 8'h01;
  filter_out_expected[1680] <= 8'h00;
  filter_out_expected[1681] <= 8'hff;
  filter_out_expected[1682] <= 8'h01;
  filter_out_expected[1683] <= 8'h01;
  filter_out_expected[1684] <= 8'hff;
  filter_out_expected[1685] <= 8'h00;
  filter_out_expected[1686] <= 8'h01;
  filter_out_expected[1687] <= 8'hff;
  filter_out_expected[1688] <= 8'h00;
  filter_out_expected[1689] <= 8'h01;
  filter_out_expected[1690] <= 8'h00;
  filter_out_expected[1691] <= 8'hff;
  filter_out_expected[1692] <= 8'h01;
  filter_out_expected[1693] <= 8'h00;
  filter_out_expected[1694] <= 8'hff;
  filter_out_expected[1695] <= 8'h01;
  filter_out_expected[1696] <= 8'h01;
  filter_out_expected[1697] <= 8'hff;
  filter_out_expected[1698] <= 8'h00;
  filter_out_expected[1699] <= 8'h01;
  filter_out_expected[1700] <= 8'hff;
  filter_out_expected[1701] <= 8'h00;
  filter_out_expected[1702] <= 8'h01;
  filter_out_expected[1703] <= 8'h00;
  filter_out_expected[1704] <= 8'hff;
  filter_out_expected[1705] <= 8'h01;
  filter_out_expected[1706] <= 8'h00;
  filter_out_expected[1707] <= 8'hff;
  filter_out_expected[1708] <= 8'h01;
  filter_out_expected[1709] <= 8'h00;
  filter_out_expected[1710] <= 8'hff;
  filter_out_expected[1711] <= 8'h01;
  filter_out_expected[1712] <= 8'h01;
  filter_out_expected[1713] <= 8'hff;
  filter_out_expected[1714] <= 8'h00;
  filter_out_expected[1715] <= 8'h01;
  filter_out_expected[1716] <= 8'hff;
  filter_out_expected[1717] <= 8'h00;
  filter_out_expected[1718] <= 8'h01;
  filter_out_expected[1719] <= 8'hff;
  filter_out_expected[1720] <= 8'hff;
  filter_out_expected[1721] <= 8'h01;
  filter_out_expected[1722] <= 8'hff;
  filter_out_expected[1723] <= 8'hff;
  filter_out_expected[1724] <= 8'h01;
  filter_out_expected[1725] <= 8'h00;
  filter_out_expected[1726] <= 8'hff;
  filter_out_expected[1727] <= 8'h01;
  filter_out_expected[1728] <= 8'h00;
  filter_out_expected[1729] <= 8'hff;
  filter_out_expected[1730] <= 8'h01;
  filter_out_expected[1731] <= 8'h00;
  filter_out_expected[1732] <= 8'hff;
  filter_out_expected[1733] <= 8'h01;
  filter_out_expected[1734] <= 8'h00;
  filter_out_expected[1735] <= 8'hff;
  filter_out_expected[1736] <= 8'h01;
  filter_out_expected[1737] <= 8'h00;
  filter_out_expected[1738] <= 8'hfe;
  filter_out_expected[1739] <= 8'h01;
  filter_out_expected[1740] <= 8'h00;
  filter_out_expected[1741] <= 8'hfe;
  filter_out_expected[1742] <= 8'h01;
  filter_out_expected[1743] <= 8'h01;
  filter_out_expected[1744] <= 8'hfe;
  filter_out_expected[1745] <= 8'h01;
  filter_out_expected[1746] <= 8'h01;
  filter_out_expected[1747] <= 8'hfe;
  filter_out_expected[1748] <= 8'h01;
  filter_out_expected[1749] <= 8'h01;
  filter_out_expected[1750] <= 8'hfe;
  filter_out_expected[1751] <= 8'h01;
  filter_out_expected[1752] <= 8'h01;
  filter_out_expected[1753] <= 8'hfe;
  filter_out_expected[1754] <= 8'h01;
  filter_out_expected[1755] <= 8'h00;
  filter_out_expected[1756] <= 8'hff;
  filter_out_expected[1757] <= 8'h01;
  filter_out_expected[1758] <= 8'h00;
  filter_out_expected[1759] <= 8'hff;
  filter_out_expected[1760] <= 8'h01;
  filter_out_expected[1761] <= 8'h00;
  filter_out_expected[1762] <= 8'hff;
  filter_out_expected[1763] <= 8'h01;
  filter_out_expected[1764] <= 8'h00;
  filter_out_expected[1765] <= 8'hff;
  filter_out_expected[1766] <= 8'h01;
  filter_out_expected[1767] <= 8'h00;
  filter_out_expected[1768] <= 8'hff;
  filter_out_expected[1769] <= 8'h01;
  filter_out_expected[1770] <= 8'hff;
  filter_out_expected[1771] <= 8'hff;
  filter_out_expected[1772] <= 8'h02;
  filter_out_expected[1773] <= 8'hff;
  filter_out_expected[1774] <= 8'h00;
  filter_out_expected[1775] <= 8'h01;
  filter_out_expected[1776] <= 8'hff;
  filter_out_expected[1777] <= 8'h00;
  filter_out_expected[1778] <= 8'h01;
  filter_out_expected[1779] <= 8'hff;
  filter_out_expected[1780] <= 8'h00;
  filter_out_expected[1781] <= 8'h01;
  filter_out_expected[1782] <= 8'hff;
  filter_out_expected[1783] <= 8'h01;
  filter_out_expected[1784] <= 8'h01;
  filter_out_expected[1785] <= 8'hff;
  filter_out_expected[1786] <= 8'h01;
  filter_out_expected[1787] <= 8'h00;
  filter_out_expected[1788] <= 8'hff;
  filter_out_expected[1789] <= 8'h01;
  filter_out_expected[1790] <= 8'h00;
  filter_out_expected[1791] <= 8'hff;
  filter_out_expected[1792] <= 8'h01;
  filter_out_expected[1793] <= 8'hff;
  filter_out_expected[1794] <= 8'h00;
  filter_out_expected[1795] <= 8'h01;
  filter_out_expected[1796] <= 8'hff;
  filter_out_expected[1797] <= 8'h00;
  filter_out_expected[1798] <= 8'h01;
  filter_out_expected[1799] <= 8'hff;
  filter_out_expected[1800] <= 8'h01;
  filter_out_expected[1801] <= 8'h00;
  filter_out_expected[1802] <= 8'hff;
  filter_out_expected[1803] <= 8'h01;
  filter_out_expected[1804] <= 8'h00;
  filter_out_expected[1805] <= 8'hff;
  filter_out_expected[1806] <= 8'h01;
  filter_out_expected[1807] <= 8'hff;
  filter_out_expected[1808] <= 8'h00;
  filter_out_expected[1809] <= 8'h01;
  filter_out_expected[1810] <= 8'hff;
  filter_out_expected[1811] <= 8'h01;
  filter_out_expected[1812] <= 8'h00;
  filter_out_expected[1813] <= 8'hff;
  filter_out_expected[1814] <= 8'h01;
  filter_out_expected[1815] <= 8'h00;
  filter_out_expected[1816] <= 8'hff;
  filter_out_expected[1817] <= 8'h01;
  filter_out_expected[1818] <= 8'hff;
  filter_out_expected[1819] <= 8'h00;
  filter_out_expected[1820] <= 8'h01;
  filter_out_expected[1821] <= 8'hff;
  filter_out_expected[1822] <= 8'h01;
  filter_out_expected[1823] <= 8'h00;
  filter_out_expected[1824] <= 8'hff;
  filter_out_expected[1825] <= 8'h01;
  filter_out_expected[1826] <= 8'hff;
  filter_out_expected[1827] <= 8'h00;
  filter_out_expected[1828] <= 8'h01;
  filter_out_expected[1829] <= 8'hff;
  filter_out_expected[1830] <= 8'h01;
  filter_out_expected[1831] <= 8'h00;
  filter_out_expected[1832] <= 8'hff;
  filter_out_expected[1833] <= 8'h01;
  filter_out_expected[1834] <= 8'hff;
  filter_out_expected[1835] <= 8'h00;
  filter_out_expected[1836] <= 8'h01;
  filter_out_expected[1837] <= 8'hff;
  filter_out_expected[1838] <= 8'h00;
  filter_out_expected[1839] <= 8'h00;
  filter_out_expected[1840] <= 8'hff;
  filter_out_expected[1841] <= 8'h01;
  filter_out_expected[1842] <= 8'hff;
  filter_out_expected[1843] <= 8'h00;
  filter_out_expected[1844] <= 8'h01;
  filter_out_expected[1845] <= 8'hff;
  filter_out_expected[1846] <= 8'h01;
  filter_out_expected[1847] <= 8'h00;
  filter_out_expected[1848] <= 8'hff;
  filter_out_expected[1849] <= 8'h01;
  filter_out_expected[1850] <= 8'hff;
  filter_out_expected[1851] <= 8'h00;
  filter_out_expected[1852] <= 8'h00;
  filter_out_expected[1853] <= 8'hff;
  filter_out_expected[1854] <= 8'h01;
  filter_out_expected[1855] <= 8'h00;
  filter_out_expected[1856] <= 8'h00;
  filter_out_expected[1857] <= 8'h01;
  filter_out_expected[1858] <= 8'hff;
  filter_out_expected[1859] <= 8'h00;
  filter_out_expected[1860] <= 8'h00;
  filter_out_expected[1861] <= 8'h00;
  filter_out_expected[1862] <= 8'h01;
  filter_out_expected[1863] <= 8'hff;
  filter_out_expected[1864] <= 8'h00;
  filter_out_expected[1865] <= 8'h00;
  filter_out_expected[1866] <= 8'hff;
  filter_out_expected[1867] <= 8'h01;
  filter_out_expected[1868] <= 8'h00;
  filter_out_expected[1869] <= 8'h00;
  filter_out_expected[1870] <= 8'h00;
  filter_out_expected[1871] <= 8'hff;
  filter_out_expected[1872] <= 8'h00;
  filter_out_expected[1873] <= 8'h00;
  filter_out_expected[1874] <= 8'h00;
  filter_out_expected[1875] <= 8'h00;
  filter_out_expected[1876] <= 8'hff;
  filter_out_expected[1877] <= 8'h00;
  filter_out_expected[1878] <= 8'h00;
  filter_out_expected[1879] <= 8'h00;
  filter_out_expected[1880] <= 8'h00;
  filter_out_expected[1881] <= 8'h00;
  filter_out_expected[1882] <= 8'h00;
  filter_out_expected[1883] <= 8'h00;
  filter_out_expected[1884] <= 8'h00;
  filter_out_expected[1885] <= 8'h00;
  filter_out_expected[1886] <= 8'h00;
  filter_out_expected[1887] <= 8'h00;
  filter_out_expected[1888] <= 8'h00;
  filter_out_expected[1889] <= 8'h00;
  filter_out_expected[1890] <= 8'h00;
  filter_out_expected[1891] <= 8'h00;
  filter_out_expected[1892] <= 8'h00;
  filter_out_expected[1893] <= 8'h00;
  filter_out_expected[1894] <= 8'h00;
  filter_out_expected[1895] <= 8'h00;
  filter_out_expected[1896] <= 8'h00;
  filter_out_expected[1897] <= 8'h00;
  filter_out_expected[1898] <= 8'h00;
  filter_out_expected[1899] <= 8'h00;
  filter_out_expected[1900] <= 8'h00;
  filter_out_expected[1901] <= 8'h00;
  filter_out_expected[1902] <= 8'h00;
  filter_out_expected[1903] <= 8'h00;
  filter_out_expected[1904] <= 8'h00;
  filter_out_expected[1905] <= 8'h00;
  filter_out_expected[1906] <= 8'h00;
  filter_out_expected[1907] <= 8'h00;
  filter_out_expected[1908] <= 8'h00;
  filter_out_expected[1909] <= 8'h00;
  filter_out_expected[1910] <= 8'h00;
  filter_out_expected[1911] <= 8'h00;
  filter_out_expected[1912] <= 8'h00;
  filter_out_expected[1913] <= 8'h00;
  filter_out_expected[1914] <= 8'h00;
  filter_out_expected[1915] <= 8'h00;
  filter_out_expected[1916] <= 8'h00;
  filter_out_expected[1917] <= 8'h00;
  filter_out_expected[1918] <= 8'h00;
  filter_out_expected[1919] <= 8'h00;
  filter_out_expected[1920] <= 8'h00;
  filter_out_expected[1921] <= 8'h00;
  filter_out_expected[1922] <= 8'h00;
  filter_out_expected[1923] <= 8'h00;
  filter_out_expected[1924] <= 8'h00;
  filter_out_expected[1925] <= 8'h00;
  filter_out_expected[1926] <= 8'h00;
  filter_out_expected[1927] <= 8'h00;
  filter_out_expected[1928] <= 8'h00;
  filter_out_expected[1929] <= 8'h00;
  filter_out_expected[1930] <= 8'h00;
  filter_out_expected[1931] <= 8'h00;
  filter_out_expected[1932] <= 8'h00;
  filter_out_expected[1933] <= 8'h00;
  filter_out_expected[1934] <= 8'h00;
  filter_out_expected[1935] <= 8'h00;
  filter_out_expected[1936] <= 8'h00;
  filter_out_expected[1937] <= 8'h00;
  filter_out_expected[1938] <= 8'h00;
  filter_out_expected[1939] <= 8'h00;
  filter_out_expected[1940] <= 8'h00;
  filter_out_expected[1941] <= 8'h00;
  filter_out_expected[1942] <= 8'h00;
  filter_out_expected[1943] <= 8'h00;
  filter_out_expected[1944] <= 8'h00;
  filter_out_expected[1945] <= 8'h00;
  filter_out_expected[1946] <= 8'h00;
  filter_out_expected[1947] <= 8'h00;
  filter_out_expected[1948] <= 8'h00;
  filter_out_expected[1949] <= 8'h00;
  filter_out_expected[1950] <= 8'hff;
  filter_out_expected[1951] <= 8'h00;
  filter_out_expected[1952] <= 8'h00;
  filter_out_expected[1953] <= 8'h00;
  filter_out_expected[1954] <= 8'h00;
  filter_out_expected[1955] <= 8'h00;
  filter_out_expected[1956] <= 8'h00;
  filter_out_expected[1957] <= 8'hff;
  filter_out_expected[1958] <= 8'h01;
  filter_out_expected[1959] <= 8'hff;
  filter_out_expected[1960] <= 8'h00;
  filter_out_expected[1961] <= 8'h00;
  filter_out_expected[1962] <= 8'h00;
  filter_out_expected[1963] <= 8'h00;
  filter_out_expected[1964] <= 8'h00;
  filter_out_expected[1965] <= 8'h01;
  filter_out_expected[1966] <= 8'hff;
  filter_out_expected[1967] <= 8'h01;
  filter_out_expected[1968] <= 8'hff;
  filter_out_expected[1969] <= 8'h00;
  filter_out_expected[1970] <= 8'h00;
  filter_out_expected[1971] <= 8'h00;
  filter_out_expected[1972] <= 8'h00;
  filter_out_expected[1973] <= 8'hff;
  filter_out_expected[1974] <= 8'h01;
  filter_out_expected[1975] <= 8'hff;
  filter_out_expected[1976] <= 8'h01;
  filter_out_expected[1977] <= 8'hff;
  filter_out_expected[1978] <= 8'h00;
  filter_out_expected[1979] <= 8'h00;
  filter_out_expected[1980] <= 8'h00;
  filter_out_expected[1981] <= 8'h01;
  filter_out_expected[1982] <= 8'hff;
  filter_out_expected[1983] <= 8'h01;
  filter_out_expected[1984] <= 8'hff;
  filter_out_expected[1985] <= 8'h01;
  filter_out_expected[1986] <= 8'hff;
  filter_out_expected[1987] <= 8'h00;
  filter_out_expected[1988] <= 8'h00;
  filter_out_expected[1989] <= 8'h00;
  filter_out_expected[1990] <= 8'h00;
  filter_out_expected[1991] <= 8'hff;
  filter_out_expected[1992] <= 8'h01;
  filter_out_expected[1993] <= 8'hff;
  filter_out_expected[1994] <= 8'h01;
  filter_out_expected[1995] <= 8'hff;
  filter_out_expected[1996] <= 8'h01;
  filter_out_expected[1997] <= 8'h00;
  filter_out_expected[1998] <= 8'h00;
  filter_out_expected[1999] <= 8'h00;
  filter_out_expected[2000] <= 8'h00;
  filter_out_expected[2001] <= 8'h01;
  filter_out_expected[2002] <= 8'hff;
  filter_out_expected[2003] <= 8'h01;
  filter_out_expected[2004] <= 8'hff;
  filter_out_expected[2005] <= 8'h01;
  filter_out_expected[2006] <= 8'hff;
  filter_out_expected[2007] <= 8'h01;
  filter_out_expected[2008] <= 8'hff;
  filter_out_expected[2009] <= 8'h00;
  filter_out_expected[2010] <= 8'h00;
  filter_out_expected[2011] <= 8'h00;
  filter_out_expected[2012] <= 8'h01;
  filter_out_expected[2013] <= 8'hff;
  filter_out_expected[2014] <= 8'h01;
  filter_out_expected[2015] <= 8'hff;
  filter_out_expected[2016] <= 8'h01;
  filter_out_expected[2017] <= 8'hff;
  filter_out_expected[2018] <= 8'h01;
  filter_out_expected[2019] <= 8'hff;
  filter_out_expected[2020] <= 8'h01;
  filter_out_expected[2021] <= 8'hff;
  filter_out_expected[2022] <= 8'h00;
  filter_out_expected[2023] <= 8'h00;
  filter_out_expected[2024] <= 8'h00;
  filter_out_expected[2025] <= 8'h00;
  filter_out_expected[2026] <= 8'hff;
  filter_out_expected[2027] <= 8'h01;
  filter_out_expected[2028] <= 8'hff;
  filter_out_expected[2029] <= 8'h01;
  filter_out_expected[2030] <= 8'hff;
  filter_out_expected[2031] <= 8'h01;
  filter_out_expected[2032] <= 8'hff;
  filter_out_expected[2033] <= 8'h01;
  filter_out_expected[2034] <= 8'hff;
  filter_out_expected[2035] <= 8'h01;
  filter_out_expected[2036] <= 8'hff;
  filter_out_expected[2037] <= 8'h01;
  filter_out_expected[2038] <= 8'h00;
  filter_out_expected[2039] <= 8'h00;
  filter_out_expected[2040] <= 8'h00;
  filter_out_expected[2041] <= 8'h00;
  filter_out_expected[2042] <= 8'h00;
  filter_out_expected[2043] <= 8'hff;
  filter_out_expected[2044] <= 8'h01;
  filter_out_expected[2045] <= 8'hff;
  filter_out_expected[2046] <= 8'h01;
  filter_out_expected[2047] <= 8'hff;
  filter_out_expected[2048] <= 8'h01;
  filter_out_expected[2049] <= 8'hff;
  filter_out_expected[2050] <= 8'h01;
  filter_out_expected[2051] <= 8'hff;
  filter_out_expected[2052] <= 8'h01;
  filter_out_expected[2053] <= 8'hff;
  filter_out_expected[2054] <= 8'h01;
  filter_out_expected[2055] <= 8'hff;
  filter_out_expected[2056] <= 8'h01;
  filter_out_expected[2057] <= 8'hff;
  filter_out_expected[2058] <= 8'h01;
  filter_out_expected[2059] <= 8'hff;
  filter_out_expected[2060] <= 8'h01;
  filter_out_expected[2061] <= 8'hff;
  filter_out_expected[2062] <= 8'h00;
  filter_out_expected[2063] <= 8'h00;
  filter_out_expected[2064] <= 8'h00;
  filter_out_expected[2065] <= 8'h00;
  filter_out_expected[2066] <= 8'h00;
  filter_out_expected[2067] <= 8'h00;
  filter_out_expected[2068] <= 8'h00;
  filter_out_expected[2069] <= 8'h01;
  filter_out_expected[2070] <= 8'hff;
  filter_out_expected[2071] <= 8'h01;
  filter_out_expected[2072] <= 8'hff;
  filter_out_expected[2073] <= 8'hff;
  filter_out_expected[2074] <= 8'hfd;
  filter_out_expected[2075] <= 8'hfe;
  filter_out_expected[2076] <= 8'hfe;
  filter_out_expected[2077] <= 8'h00;
  filter_out_expected[2078] <= 8'hfe;
  filter_out_expected[2079] <= 8'hfd;
  filter_out_expected[2080] <= 8'hfb;
  filter_out_expected[2081] <= 8'hfc;
  filter_out_expected[2082] <= 8'h00;
  filter_out_expected[2083] <= 8'h01;
  filter_out_expected[2084] <= 8'h02;
  filter_out_expected[2085] <= 8'h04;
  filter_out_expected[2086] <= 8'h05;
  filter_out_expected[2087] <= 8'h04;
  filter_out_expected[2088] <= 8'h03;
  filter_out_expected[2089] <= 8'h01;
  filter_out_expected[2090] <= 8'h03;
  filter_out_expected[2091] <= 8'h08;
  filter_out_expected[2092] <= 8'h09;
  filter_out_expected[2093] <= 8'h06;
  filter_out_expected[2094] <= 8'h05;
  filter_out_expected[2095] <= 8'h05;
  filter_out_expected[2096] <= 8'h08;
  filter_out_expected[2097] <= 8'h09;
  filter_out_expected[2098] <= 8'h07;
  filter_out_expected[2099] <= 8'h03;
  filter_out_expected[2100] <= 8'h05;
  filter_out_expected[2101] <= 8'h05;
  filter_out_expected[2102] <= 8'h04;
  filter_out_expected[2103] <= 8'h00;
  filter_out_expected[2104] <= 8'hfc;
  filter_out_expected[2105] <= 8'hfb;
  filter_out_expected[2106] <= 8'h01;
  filter_out_expected[2107] <= 8'h06;
  filter_out_expected[2108] <= 8'h09;
  filter_out_expected[2109] <= 8'h07;
  filter_out_expected[2110] <= 8'h02;
  filter_out_expected[2111] <= 8'hfe;
  filter_out_expected[2112] <= 8'hfc;
  filter_out_expected[2113] <= 8'hfd;
  filter_out_expected[2114] <= 8'hff;
  filter_out_expected[2115] <= 8'hfe;
  filter_out_expected[2116] <= 8'hfd;
  filter_out_expected[2117] <= 8'hfa;
  filter_out_expected[2118] <= 8'hfb;
  filter_out_expected[2119] <= 8'h03;
  filter_out_expected[2120] <= 8'h06;
  filter_out_expected[2121] <= 8'h04;
  filter_out_expected[2122] <= 8'h01;
  filter_out_expected[2123] <= 8'hfd;
  filter_out_expected[2124] <= 8'hff;
  filter_out_expected[2125] <= 8'h08;
  filter_out_expected[2126] <= 8'h0e;
  filter_out_expected[2127] <= 8'h10;
  filter_out_expected[2128] <= 8'h0f;
  filter_out_expected[2129] <= 8'h0a;
  filter_out_expected[2130] <= 8'h08;
  filter_out_expected[2131] <= 8'h09;
  filter_out_expected[2132] <= 8'h0c;
  filter_out_expected[2133] <= 8'h0e;
  filter_out_expected[2134] <= 8'h0d;
  filter_out_expected[2135] <= 8'h0a;
  filter_out_expected[2136] <= 8'h09;
  filter_out_expected[2137] <= 8'h06;
  filter_out_expected[2138] <= 8'h03;
  filter_out_expected[2139] <= 8'h03;
  filter_out_expected[2140] <= 8'h02;
  filter_out_expected[2141] <= 8'h04;
  filter_out_expected[2142] <= 8'h08;
  filter_out_expected[2143] <= 8'h0c;
  filter_out_expected[2144] <= 8'h0e;
  filter_out_expected[2145] <= 8'h0d;
  filter_out_expected[2146] <= 8'h03;
  filter_out_expected[2147] <= 8'hfa;
  filter_out_expected[2148] <= 8'hf7;
  filter_out_expected[2149] <= 8'hfd;
  filter_out_expected[2150] <= 8'h07;
  filter_out_expected[2151] <= 8'h0d;
  filter_out_expected[2152] <= 8'h0c;
  filter_out_expected[2153] <= 8'h07;
  filter_out_expected[2154] <= 8'h04;
  filter_out_expected[2155] <= 8'h04;
  filter_out_expected[2156] <= 8'h02;
  filter_out_expected[2157] <= 8'h00;
  filter_out_expected[2158] <= 8'hff;
  filter_out_expected[2159] <= 8'hfb;
  filter_out_expected[2160] <= 8'hfd;
  filter_out_expected[2161] <= 8'hfe;
  filter_out_expected[2162] <= 8'hfd;
  filter_out_expected[2163] <= 8'hfa;
  filter_out_expected[2164] <= 8'hf6;
  filter_out_expected[2165] <= 8'hf2;
  filter_out_expected[2166] <= 8'hf4;
  filter_out_expected[2167] <= 8'hf6;
  filter_out_expected[2168] <= 8'hf7;
  filter_out_expected[2169] <= 8'hf6;
  filter_out_expected[2170] <= 8'hf8;
  filter_out_expected[2171] <= 8'hfc;
  filter_out_expected[2172] <= 8'h03;
  filter_out_expected[2173] <= 8'h06;
  filter_out_expected[2174] <= 8'h09;
  filter_out_expected[2175] <= 8'h05;
  filter_out_expected[2176] <= 8'h05;
  filter_out_expected[2177] <= 8'h06;
  filter_out_expected[2178] <= 8'h06;
  filter_out_expected[2179] <= 8'h03;
  filter_out_expected[2180] <= 8'hff;
  filter_out_expected[2181] <= 8'hfb;
  filter_out_expected[2182] <= 8'hfa;
  filter_out_expected[2183] <= 8'hfd;
  filter_out_expected[2184] <= 8'hfe;
  filter_out_expected[2185] <= 8'h01;
  filter_out_expected[2186] <= 8'h02;
  filter_out_expected[2187] <= 8'h00;
  filter_out_expected[2188] <= 8'hfc;
  filter_out_expected[2189] <= 8'hf9;
  filter_out_expected[2190] <= 8'hf7;
  filter_out_expected[2191] <= 8'hf7;
  filter_out_expected[2192] <= 8'hf8;
  filter_out_expected[2193] <= 8'hfa;
  filter_out_expected[2194] <= 8'hff;
  filter_out_expected[2195] <= 8'h05;
  filter_out_expected[2196] <= 8'h0a;
  filter_out_expected[2197] <= 8'h09;
  filter_out_expected[2198] <= 8'h03;
  filter_out_expected[2199] <= 8'hfb;
  filter_out_expected[2200] <= 8'hfb;
  filter_out_expected[2201] <= 8'h01;
  filter_out_expected[2202] <= 8'h08;
  filter_out_expected[2203] <= 8'h08;
  filter_out_expected[2204] <= 8'h01;
  filter_out_expected[2205] <= 8'hfb;
  filter_out_expected[2206] <= 8'hfa;
  filter_out_expected[2207] <= 8'hfc;
  filter_out_expected[2208] <= 8'hfc;
  filter_out_expected[2209] <= 8'hfa;
  filter_out_expected[2210] <= 8'hf9;
  filter_out_expected[2211] <= 8'hfa;
  filter_out_expected[2212] <= 8'h00;
  filter_out_expected[2213] <= 8'h01;
  filter_out_expected[2214] <= 8'h03;
  filter_out_expected[2215] <= 8'h02;
  filter_out_expected[2216] <= 8'h04;
  filter_out_expected[2217] <= 8'h04;
  filter_out_expected[2218] <= 8'h07;
  filter_out_expected[2219] <= 8'h04;
  filter_out_expected[2220] <= 8'h03;
  filter_out_expected[2221] <= 8'hff;
  filter_out_expected[2222] <= 8'hfb;
  filter_out_expected[2223] <= 8'hf6;
  filter_out_expected[2224] <= 8'hf8;
  filter_out_expected[2225] <= 8'hf8;
  filter_out_expected[2226] <= 8'hfd;
  filter_out_expected[2227] <= 8'hfe;
  filter_out_expected[2228] <= 8'h01;
  filter_out_expected[2229] <= 8'h04;
  filter_out_expected[2230] <= 8'h06;
  filter_out_expected[2231] <= 8'h05;
  filter_out_expected[2232] <= 8'h03;
  filter_out_expected[2233] <= 8'h03;
  filter_out_expected[2234] <= 8'h02;
  filter_out_expected[2235] <= 8'h02;
  filter_out_expected[2236] <= 8'h00;
  filter_out_expected[2237] <= 8'h04;
  filter_out_expected[2238] <= 8'h07;
  filter_out_expected[2239] <= 8'h06;
  filter_out_expected[2240] <= 8'hfe;
  filter_out_expected[2241] <= 8'hf7;
  filter_out_expected[2242] <= 8'hf7;
  filter_out_expected[2243] <= 8'hff;
  filter_out_expected[2244] <= 8'h05;
  filter_out_expected[2245] <= 8'h08;
  filter_out_expected[2246] <= 8'h07;
  filter_out_expected[2247] <= 8'h09;
  filter_out_expected[2248] <= 8'h08;
  filter_out_expected[2249] <= 8'h03;
  filter_out_expected[2250] <= 8'hfd;
  filter_out_expected[2251] <= 8'hff;
  filter_out_expected[2252] <= 8'h05;
  filter_out_expected[2253] <= 8'h0a;
  filter_out_expected[2254] <= 8'h06;
  filter_out_expected[2255] <= 8'h01;
  filter_out_expected[2256] <= 8'h00;
  filter_out_expected[2257] <= 8'h02;
  filter_out_expected[2258] <= 8'h02;
  filter_out_expected[2259] <= 8'hfe;
  filter_out_expected[2260] <= 8'hfb;
  filter_out_expected[2261] <= 8'hfe;
  filter_out_expected[2262] <= 8'h05;
  filter_out_expected[2263] <= 8'h09;
  filter_out_expected[2264] <= 8'h07;
  filter_out_expected[2265] <= 8'h02;
  filter_out_expected[2266] <= 8'h02;
  filter_out_expected[2267] <= 8'h04;
  filter_out_expected[2268] <= 8'h05;
  filter_out_expected[2269] <= 8'h03;
  filter_out_expected[2270] <= 8'hfe;
  filter_out_expected[2271] <= 8'hfd;
  filter_out_expected[2272] <= 8'h00;
  filter_out_expected[2273] <= 8'h07;
  filter_out_expected[2274] <= 8'h0d;
  filter_out_expected[2275] <= 8'h0e;
  filter_out_expected[2276] <= 8'h09;
  filter_out_expected[2277] <= 8'h02;
  filter_out_expected[2278] <= 8'hfb;
  filter_out_expected[2279] <= 8'hf5;
  filter_out_expected[2280] <= 8'hf1;
  filter_out_expected[2281] <= 8'hf1;
  filter_out_expected[2282] <= 8'hf3;
  filter_out_expected[2283] <= 8'hf8;
  filter_out_expected[2284] <= 8'hfe;
  filter_out_expected[2285] <= 8'h06;
  filter_out_expected[2286] <= 8'h0a;
  filter_out_expected[2287] <= 8'h0c;
  filter_out_expected[2288] <= 8'h0b;
  filter_out_expected[2289] <= 8'h0a;
  filter_out_expected[2290] <= 8'h07;
  filter_out_expected[2291] <= 8'h07;
  filter_out_expected[2292] <= 8'h02;
  filter_out_expected[2293] <= 8'hfe;
  filter_out_expected[2294] <= 8'hfe;
  filter_out_expected[2295] <= 8'h00;
  filter_out_expected[2296] <= 8'hff;
  filter_out_expected[2297] <= 8'hfe;
  filter_out_expected[2298] <= 8'hfc;
  filter_out_expected[2299] <= 8'hfa;
  filter_out_expected[2300] <= 8'hfb;
  filter_out_expected[2301] <= 8'hfe;
  filter_out_expected[2302] <= 8'h00;
  filter_out_expected[2303] <= 8'h03;
  filter_out_expected[2304] <= 8'h06;
  filter_out_expected[2305] <= 8'h06;
  filter_out_expected[2306] <= 8'h02;
  filter_out_expected[2307] <= 8'hff;
  filter_out_expected[2308] <= 8'hf9;
  filter_out_expected[2309] <= 8'hf8;
  filter_out_expected[2310] <= 8'hf9;
  filter_out_expected[2311] <= 8'h00;
  filter_out_expected[2312] <= 8'h01;
  filter_out_expected[2313] <= 8'h03;
  filter_out_expected[2314] <= 8'h03;
  filter_out_expected[2315] <= 8'h03;
  filter_out_expected[2316] <= 8'hfe;
  filter_out_expected[2317] <= 8'hf7;
  filter_out_expected[2318] <= 8'hf2;
  filter_out_expected[2319] <= 8'hf3;
  filter_out_expected[2320] <= 8'hf9;
  filter_out_expected[2321] <= 8'hfe;
  filter_out_expected[2322] <= 8'h01;
  filter_out_expected[2323] <= 8'hff;
  filter_out_expected[2324] <= 8'hfb;
  filter_out_expected[2325] <= 8'hf5;
  filter_out_expected[2326] <= 8'hf2;
  filter_out_expected[2327] <= 8'hf4;
  filter_out_expected[2328] <= 8'hf7;
  filter_out_expected[2329] <= 8'hf6;
  filter_out_expected[2330] <= 8'hf3;
  filter_out_expected[2331] <= 8'hf4;
  filter_out_expected[2332] <= 8'hfb;
  filter_out_expected[2333] <= 8'h03;
  filter_out_expected[2334] <= 8'h09;
  filter_out_expected[2335] <= 8'h0a;
  filter_out_expected[2336] <= 8'h06;
  filter_out_expected[2337] <= 8'h02;
  filter_out_expected[2338] <= 8'hfe;
  filter_out_expected[2339] <= 8'hfa;
  filter_out_expected[2340] <= 8'hf4;
  filter_out_expected[2341] <= 8'hf4;
  filter_out_expected[2342] <= 8'hfb;
  filter_out_expected[2343] <= 8'h03;
  filter_out_expected[2344] <= 8'h05;
  filter_out_expected[2345] <= 8'h03;
  filter_out_expected[2346] <= 8'hfe;
  filter_out_expected[2347] <= 8'hff;
  filter_out_expected[2348] <= 8'h02;
  filter_out_expected[2349] <= 8'h03;
  filter_out_expected[2350] <= 8'h00;
  filter_out_expected[2351] <= 8'h00;
  filter_out_expected[2352] <= 8'h01;
  filter_out_expected[2353] <= 8'h07;
  filter_out_expected[2354] <= 8'h0a;
  filter_out_expected[2355] <= 8'h0b;
  filter_out_expected[2356] <= 8'h08;
  filter_out_expected[2357] <= 8'h04;
  filter_out_expected[2358] <= 8'h04;
  filter_out_expected[2359] <= 8'h04;
  filter_out_expected[2360] <= 8'h01;
  filter_out_expected[2361] <= 8'h02;
  filter_out_expected[2362] <= 8'hff;
  filter_out_expected[2363] <= 8'hfc;
  filter_out_expected[2364] <= 8'hfb;
  filter_out_expected[2365] <= 8'hfa;
  filter_out_expected[2366] <= 8'hfa;
  filter_out_expected[2367] <= 8'hff;
  filter_out_expected[2368] <= 8'h03;
  filter_out_expected[2369] <= 8'h05;
  filter_out_expected[2370] <= 8'h08;
  filter_out_expected[2371] <= 8'h06;
  filter_out_expected[2372] <= 8'h04;
  filter_out_expected[2373] <= 8'hff;
  filter_out_expected[2374] <= 8'hfc;
  filter_out_expected[2375] <= 8'hfc;
  filter_out_expected[2376] <= 8'h03;
  filter_out_expected[2377] <= 8'h08;
  filter_out_expected[2378] <= 8'h09;
  filter_out_expected[2379] <= 8'h05;
  filter_out_expected[2380] <= 8'h04;
  filter_out_expected[2381] <= 8'h05;
  filter_out_expected[2382] <= 8'h0a;
  filter_out_expected[2383] <= 8'h0a;
  filter_out_expected[2384] <= 8'h04;
  filter_out_expected[2385] <= 8'hfb;
  filter_out_expected[2386] <= 8'hf6;
  filter_out_expected[2387] <= 8'hf5;
  filter_out_expected[2388] <= 8'hf7;
  filter_out_expected[2389] <= 8'hfb;
  filter_out_expected[2390] <= 8'hfb;
  filter_out_expected[2391] <= 8'hfb;
  filter_out_expected[2392] <= 8'hf9;
  filter_out_expected[2393] <= 8'hf7;
  filter_out_expected[2394] <= 8'hf4;
  filter_out_expected[2395] <= 8'hf6;
  filter_out_expected[2396] <= 8'hf6;
  filter_out_expected[2397] <= 8'hf7;
  filter_out_expected[2398] <= 8'hf4;
  filter_out_expected[2399] <= 8'hf1;
  filter_out_expected[2400] <= 8'hf1;
  filter_out_expected[2401] <= 8'hf7;
  filter_out_expected[2402] <= 8'hfd;
  filter_out_expected[2403] <= 8'h02;
  filter_out_expected[2404] <= 8'h01;
  filter_out_expected[2405] <= 8'h00;
  filter_out_expected[2406] <= 8'h02;
  filter_out_expected[2407] <= 8'h09;
  filter_out_expected[2408] <= 8'h09;
  filter_out_expected[2409] <= 8'h08;
  filter_out_expected[2410] <= 8'h01;
  filter_out_expected[2411] <= 8'hfb;
  filter_out_expected[2412] <= 8'hf9;
  filter_out_expected[2413] <= 8'hfb;
  filter_out_expected[2414] <= 8'hfc;
  filter_out_expected[2415] <= 8'hfd;
  filter_out_expected[2416] <= 8'h01;
  filter_out_expected[2417] <= 8'h03;
  filter_out_expected[2418] <= 8'h07;
  filter_out_expected[2419] <= 8'h08;
  filter_out_expected[2420] <= 8'h02;
  filter_out_expected[2421] <= 8'hfa;
  filter_out_expected[2422] <= 8'hf8;
  filter_out_expected[2423] <= 8'hf9;
  filter_out_expected[2424] <= 8'hfb;
  filter_out_expected[2425] <= 8'hfb;
  filter_out_expected[2426] <= 8'hf9;
  filter_out_expected[2427] <= 8'hfa;
  filter_out_expected[2428] <= 8'hff;
  filter_out_expected[2429] <= 8'h04;
  filter_out_expected[2430] <= 8'h08;
  filter_out_expected[2431] <= 8'h08;
  filter_out_expected[2432] <= 8'h03;
  filter_out_expected[2433] <= 8'hfe;
  filter_out_expected[2434] <= 8'hfd;
  filter_out_expected[2435] <= 8'hfd;
  filter_out_expected[2436] <= 8'h00;
  filter_out_expected[2437] <= 8'h01;
  filter_out_expected[2438] <= 8'h01;
  filter_out_expected[2439] <= 8'h03;
  filter_out_expected[2440] <= 8'h06;
  filter_out_expected[2441] <= 8'h08;
  filter_out_expected[2442] <= 8'h09;
  filter_out_expected[2443] <= 8'h05;
  filter_out_expected[2444] <= 8'h01;
  filter_out_expected[2445] <= 8'hfc;
  filter_out_expected[2446] <= 8'hfe;
  filter_out_expected[2447] <= 8'h01;
  filter_out_expected[2448] <= 8'h05;
  filter_out_expected[2449] <= 8'h03;
  filter_out_expected[2450] <= 8'hff;
  filter_out_expected[2451] <= 8'hfc;
  filter_out_expected[2452] <= 8'hfa;
  filter_out_expected[2453] <= 8'hfb;
  filter_out_expected[2454] <= 8'hff;
  filter_out_expected[2455] <= 8'h02;
  filter_out_expected[2456] <= 8'h02;
  filter_out_expected[2457] <= 8'h04;
  filter_out_expected[2458] <= 8'h04;
  filter_out_expected[2459] <= 8'h04;
  filter_out_expected[2460] <= 8'h01;
  filter_out_expected[2461] <= 8'hfc;
  filter_out_expected[2462] <= 8'hf6;
  filter_out_expected[2463] <= 8'hf9;
  filter_out_expected[2464] <= 8'hfc;
  filter_out_expected[2465] <= 8'hfe;
  filter_out_expected[2466] <= 8'hfd;
  filter_out_expected[2467] <= 8'hfd;
  filter_out_expected[2468] <= 8'hfb;
  filter_out_expected[2469] <= 8'hff;
  filter_out_expected[2470] <= 8'hff;
  filter_out_expected[2471] <= 8'hfd;
  filter_out_expected[2472] <= 8'hf9;
  filter_out_expected[2473] <= 8'hf8;
  filter_out_expected[2474] <= 8'hfa;
  filter_out_expected[2475] <= 8'hff;
  filter_out_expected[2476] <= 8'h01;
  filter_out_expected[2477] <= 8'h02;
  filter_out_expected[2478] <= 8'h03;
  filter_out_expected[2479] <= 8'h06;
  filter_out_expected[2480] <= 8'h0a;
  filter_out_expected[2481] <= 8'h0a;
  filter_out_expected[2482] <= 8'h07;
  filter_out_expected[2483] <= 8'h02;
  filter_out_expected[2484] <= 8'hfe;
  filter_out_expected[2485] <= 8'hfd;
  filter_out_expected[2486] <= 8'h00;
  filter_out_expected[2487] <= 8'h02;
  filter_out_expected[2488] <= 8'h00;
  filter_out_expected[2489] <= 8'hff;
  filter_out_expected[2490] <= 8'hfe;
  filter_out_expected[2491] <= 8'hfe;
  filter_out_expected[2492] <= 8'hff;
  filter_out_expected[2493] <= 8'h00;
  filter_out_expected[2494] <= 8'h01;
  filter_out_expected[2495] <= 8'h00;
  filter_out_expected[2496] <= 8'hfc;
  filter_out_expected[2497] <= 8'hf8;
  filter_out_expected[2498] <= 8'hf7;
  filter_out_expected[2499] <= 8'hfc;
  filter_out_expected[2500] <= 8'hfe;
  filter_out_expected[2501] <= 8'h00;
  filter_out_expected[2502] <= 8'h01;
  filter_out_expected[2503] <= 8'h02;
  filter_out_expected[2504] <= 8'h02;
  filter_out_expected[2505] <= 8'h01;
  filter_out_expected[2506] <= 8'hff;
  filter_out_expected[2507] <= 8'hff;
  filter_out_expected[2508] <= 8'hff;
  filter_out_expected[2509] <= 8'hf9;
  filter_out_expected[2510] <= 8'hf8;
  filter_out_expected[2511] <= 8'hfa;
  filter_out_expected[2512] <= 8'hff;
  filter_out_expected[2513] <= 8'h01;
  filter_out_expected[2514] <= 8'hff;
  filter_out_expected[2515] <= 8'hf9;
  filter_out_expected[2516] <= 8'hf9;
  filter_out_expected[2517] <= 8'hfc;
  filter_out_expected[2518] <= 8'hff;
  filter_out_expected[2519] <= 8'h01;
  filter_out_expected[2520] <= 8'h05;
  filter_out_expected[2521] <= 8'h09;
  filter_out_expected[2522] <= 8'h0a;
  filter_out_expected[2523] <= 8'h04;
  filter_out_expected[2524] <= 8'hfd;
  filter_out_expected[2525] <= 8'hfc;
  filter_out_expected[2526] <= 8'h01;
  filter_out_expected[2527] <= 8'h07;
  filter_out_expected[2528] <= 8'h08;
  filter_out_expected[2529] <= 8'h04;
  filter_out_expected[2530] <= 8'h04;
  filter_out_expected[2531] <= 8'h06;
  filter_out_expected[2532] <= 8'h09;
  filter_out_expected[2533] <= 8'h07;
  filter_out_expected[2534] <= 8'h03;
  filter_out_expected[2535] <= 8'h00;
  filter_out_expected[2536] <= 8'h00;
  filter_out_expected[2537] <= 8'h03;
  filter_out_expected[2538] <= 8'h08;
  filter_out_expected[2539] <= 8'h0d;
  filter_out_expected[2540] <= 8'h12;
  filter_out_expected[2541] <= 8'h14;
  filter_out_expected[2542] <= 8'h0e;
  filter_out_expected[2543] <= 8'h03;
  filter_out_expected[2544] <= 8'hf6;
  filter_out_expected[2545] <= 8'hee;
  filter_out_expected[2546] <= 8'heb;
  filter_out_expected[2547] <= 8'hee;
  filter_out_expected[2548] <= 8'hf1;
  filter_out_expected[2549] <= 8'hf6;
  filter_out_expected[2550] <= 8'hfd;
  filter_out_expected[2551] <= 8'h02;
  filter_out_expected[2552] <= 8'h03;
  filter_out_expected[2553] <= 8'h03;
  filter_out_expected[2554] <= 8'h01;
  filter_out_expected[2555] <= 8'hfe;
  filter_out_expected[2556] <= 8'hfd;
  filter_out_expected[2557] <= 8'hfd;
  filter_out_expected[2558] <= 8'hfe;
  filter_out_expected[2559] <= 8'h03;
  filter_out_expected[2560] <= 8'h06;
  filter_out_expected[2561] <= 8'h05;
  filter_out_expected[2562] <= 8'h03;
  filter_out_expected[2563] <= 8'h04;
  filter_out_expected[2564] <= 8'h03;
  filter_out_expected[2565] <= 8'h00;
  filter_out_expected[2566] <= 8'hfc;
  filter_out_expected[2567] <= 8'hfa;
  filter_out_expected[2568] <= 8'hfd;
  filter_out_expected[2569] <= 8'h04;
  filter_out_expected[2570] <= 8'h06;
  filter_out_expected[2571] <= 8'h05;
  filter_out_expected[2572] <= 8'h04;
  filter_out_expected[2573] <= 8'h05;
  filter_out_expected[2574] <= 8'h06;
  filter_out_expected[2575] <= 8'h06;
  filter_out_expected[2576] <= 8'h04;
  filter_out_expected[2577] <= 8'h00;
  filter_out_expected[2578] <= 8'hfa;
  filter_out_expected[2579] <= 8'hf4;
  filter_out_expected[2580] <= 8'hf3;
  filter_out_expected[2581] <= 8'hf6;
  filter_out_expected[2582] <= 8'hfd;
  filter_out_expected[2583] <= 8'h04;
  filter_out_expected[2584] <= 8'h09;
  filter_out_expected[2585] <= 8'h0d;
  filter_out_expected[2586] <= 8'h0e;
  filter_out_expected[2587] <= 8'h07;
  filter_out_expected[2588] <= 8'h04;
  filter_out_expected[2589] <= 8'h03;
  filter_out_expected[2590] <= 8'h08;
  filter_out_expected[2591] <= 8'h0c;
  filter_out_expected[2592] <= 8'h07;
  filter_out_expected[2593] <= 8'h00;
  filter_out_expected[2594] <= 8'hfb;
  filter_out_expected[2595] <= 8'hf9;
  filter_out_expected[2596] <= 8'hfc;
  filter_out_expected[2597] <= 8'h01;
  filter_out_expected[2598] <= 8'h04;
  filter_out_expected[2599] <= 8'h05;
  filter_out_expected[2600] <= 8'h02;
  filter_out_expected[2601] <= 8'hfd;
  filter_out_expected[2602] <= 8'hf8;
  filter_out_expected[2603] <= 8'hf6;
  filter_out_expected[2604] <= 8'hfa;
  filter_out_expected[2605] <= 8'hfe;
  filter_out_expected[2606] <= 8'hfe;
  filter_out_expected[2607] <= 8'hfd;
  filter_out_expected[2608] <= 8'hfa;
  filter_out_expected[2609] <= 8'hf8;
  filter_out_expected[2610] <= 8'hfa;
  filter_out_expected[2611] <= 8'hf9;
  filter_out_expected[2612] <= 8'hfb;
  filter_out_expected[2613] <= 8'hfe;
  filter_out_expected[2614] <= 8'hfd;
  filter_out_expected[2615] <= 8'hfb;
  filter_out_expected[2616] <= 8'hfd;
  filter_out_expected[2617] <= 8'hff;
  filter_out_expected[2618] <= 8'h04;
  filter_out_expected[2619] <= 8'h06;
  filter_out_expected[2620] <= 8'h02;
  filter_out_expected[2621] <= 8'hff;
  filter_out_expected[2622] <= 8'hfc;
  filter_out_expected[2623] <= 8'hfd;
  filter_out_expected[2624] <= 8'h01;
  filter_out_expected[2625] <= 8'h03;
  filter_out_expected[2626] <= 8'h04;
  filter_out_expected[2627] <= 8'h02;
  filter_out_expected[2628] <= 8'h01;
  filter_out_expected[2629] <= 8'h02;
  filter_out_expected[2630] <= 8'h04;
  filter_out_expected[2631] <= 8'h01;
  filter_out_expected[2632] <= 8'h03;
  filter_out_expected[2633] <= 8'h02;
  filter_out_expected[2634] <= 8'h04;
  filter_out_expected[2635] <= 8'h07;
  filter_out_expected[2636] <= 8'h08;
  filter_out_expected[2637] <= 8'h09;
  filter_out_expected[2638] <= 8'h08;
  filter_out_expected[2639] <= 8'h02;
  filter_out_expected[2640] <= 8'hfd;
  filter_out_expected[2641] <= 8'hfb;
  filter_out_expected[2642] <= 8'h00;
  filter_out_expected[2643] <= 8'h08;
  filter_out_expected[2644] <= 8'h0b;
  filter_out_expected[2645] <= 8'h09;
  filter_out_expected[2646] <= 8'h03;
  filter_out_expected[2647] <= 8'hff;
  filter_out_expected[2648] <= 8'hff;
  filter_out_expected[2649] <= 8'h03;
  filter_out_expected[2650] <= 8'h04;
  filter_out_expected[2651] <= 8'h04;
  filter_out_expected[2652] <= 8'hff;
  filter_out_expected[2653] <= 8'hff;
  filter_out_expected[2654] <= 8'h02;
  filter_out_expected[2655] <= 8'h07;
  filter_out_expected[2656] <= 8'h06;
  filter_out_expected[2657] <= 8'h01;
  filter_out_expected[2658] <= 8'hfa;
  filter_out_expected[2659] <= 8'hfb;
  filter_out_expected[2660] <= 8'hfe;
  filter_out_expected[2661] <= 8'h02;
  filter_out_expected[2662] <= 8'h04;
  filter_out_expected[2663] <= 8'h05;
  filter_out_expected[2664] <= 8'h06;
  filter_out_expected[2665] <= 8'h05;
  filter_out_expected[2666] <= 8'hff;
  filter_out_expected[2667] <= 8'hfd;
  filter_out_expected[2668] <= 8'hff;
  filter_out_expected[2669] <= 8'h01;
  filter_out_expected[2670] <= 8'h03;
  filter_out_expected[2671] <= 8'h02;
  filter_out_expected[2672] <= 8'hfc;
  filter_out_expected[2673] <= 8'hf7;
  filter_out_expected[2674] <= 8'hf4;
  filter_out_expected[2675] <= 8'hf2;
  filter_out_expected[2676] <= 8'hf4;
  filter_out_expected[2677] <= 8'hf6;
  filter_out_expected[2678] <= 8'hf6;
  filter_out_expected[2679] <= 8'hf5;
  filter_out_expected[2680] <= 8'hf7;
  filter_out_expected[2681] <= 8'hfa;
  filter_out_expected[2682] <= 8'hfd;
  filter_out_expected[2683] <= 8'hff;
  filter_out_expected[2684] <= 8'hff;
  filter_out_expected[2685] <= 8'hfd;
  filter_out_expected[2686] <= 8'hf9;
  filter_out_expected[2687] <= 8'hf7;
  filter_out_expected[2688] <= 8'hf7;
  filter_out_expected[2689] <= 8'hfa;
  filter_out_expected[2690] <= 8'hff;
  filter_out_expected[2691] <= 8'h06;
  filter_out_expected[2692] <= 8'h0a;
  filter_out_expected[2693] <= 8'h0e;
  filter_out_expected[2694] <= 8'h0f;
  filter_out_expected[2695] <= 8'h0e;
  filter_out_expected[2696] <= 8'h0f;
  filter_out_expected[2697] <= 8'h0b;
  filter_out_expected[2698] <= 8'h03;
  filter_out_expected[2699] <= 8'h00;
  filter_out_expected[2700] <= 8'h01;
  filter_out_expected[2701] <= 8'h05;
  filter_out_expected[2702] <= 8'h09;
  filter_out_expected[2703] <= 8'h08;
  filter_out_expected[2704] <= 8'h02;
  filter_out_expected[2705] <= 8'hfe;
  filter_out_expected[2706] <= 8'hfa;
  filter_out_expected[2707] <= 8'hf5;
  filter_out_expected[2708] <= 8'hf4;
  filter_out_expected[2709] <= 8'hf4;
  filter_out_expected[2710] <= 8'hfa;
  filter_out_expected[2711] <= 8'h00;
  filter_out_expected[2712] <= 8'h08;
  filter_out_expected[2713] <= 8'h09;
  filter_out_expected[2714] <= 8'h07;
  filter_out_expected[2715] <= 8'h05;
  filter_out_expected[2716] <= 8'h07;
  filter_out_expected[2717] <= 8'h0a;
  filter_out_expected[2718] <= 8'h0e;
  filter_out_expected[2719] <= 8'h0f;
  filter_out_expected[2720] <= 8'h0d;
  filter_out_expected[2721] <= 8'h0d;
  filter_out_expected[2722] <= 8'h0e;
  filter_out_expected[2723] <= 8'h10;
  filter_out_expected[2724] <= 8'h12;
  filter_out_expected[2725] <= 8'h0f;
  filter_out_expected[2726] <= 8'h08;
  filter_out_expected[2727] <= 8'h05;
  filter_out_expected[2728] <= 8'h01;
  filter_out_expected[2729] <= 8'hfd;
  filter_out_expected[2730] <= 8'hf9;
  filter_out_expected[2731] <= 8'hf7;
  filter_out_expected[2732] <= 8'hf6;
  filter_out_expected[2733] <= 8'hfa;
  filter_out_expected[2734] <= 8'hfe;
  filter_out_expected[2735] <= 8'h00;
  filter_out_expected[2736] <= 8'h00;
  filter_out_expected[2737] <= 8'hfe;
  filter_out_expected[2738] <= 8'hfd;
  filter_out_expected[2739] <= 8'h00;
  filter_out_expected[2740] <= 8'h04;
  filter_out_expected[2741] <= 8'h01;
  filter_out_expected[2742] <= 8'hfc;
  filter_out_expected[2743] <= 8'hfb;
  filter_out_expected[2744] <= 8'h01;
  filter_out_expected[2745] <= 8'h09;
  filter_out_expected[2746] <= 8'h0c;
  filter_out_expected[2747] <= 8'h08;
  filter_out_expected[2748] <= 8'h04;
  filter_out_expected[2749] <= 8'h01;
  filter_out_expected[2750] <= 8'h02;
  filter_out_expected[2751] <= 8'h06;
  filter_out_expected[2752] <= 8'h06;
  filter_out_expected[2753] <= 8'h02;
  filter_out_expected[2754] <= 8'hfd;
  filter_out_expected[2755] <= 8'hfa;
  filter_out_expected[2756] <= 8'hfd;
  filter_out_expected[2757] <= 8'h01;
  filter_out_expected[2758] <= 8'h02;
  filter_out_expected[2759] <= 8'hfe;
  filter_out_expected[2760] <= 8'hf8;
  filter_out_expected[2761] <= 8'hf8;
  filter_out_expected[2762] <= 8'hfb;
  filter_out_expected[2763] <= 8'hff;
  filter_out_expected[2764] <= 8'h03;
  filter_out_expected[2765] <= 8'h02;
  filter_out_expected[2766] <= 8'hfe;
  filter_out_expected[2767] <= 8'hfd;
  filter_out_expected[2768] <= 8'hfe;
  filter_out_expected[2769] <= 8'hfe;
  filter_out_expected[2770] <= 8'hff;
  filter_out_expected[2771] <= 8'h01;
  filter_out_expected[2772] <= 8'h05;
  filter_out_expected[2773] <= 8'h06;
  filter_out_expected[2774] <= 8'h03;
  filter_out_expected[2775] <= 8'hfc;
  filter_out_expected[2776] <= 8'hfa;
  filter_out_expected[2777] <= 8'hfd;
  filter_out_expected[2778] <= 8'h00;
  filter_out_expected[2779] <= 8'h00;
  filter_out_expected[2780] <= 8'hfe;
  filter_out_expected[2781] <= 8'h00;
  filter_out_expected[2782] <= 8'h07;
  filter_out_expected[2783] <= 8'h0e;
  filter_out_expected[2784] <= 8'h10;
  filter_out_expected[2785] <= 8'h10;
  filter_out_expected[2786] <= 8'h0f;
  filter_out_expected[2787] <= 8'h0a;
  filter_out_expected[2788] <= 8'h04;
  filter_out_expected[2789] <= 8'hfb;
  filter_out_expected[2790] <= 8'hf7;
  filter_out_expected[2791] <= 8'hf8;
  filter_out_expected[2792] <= 8'hfd;
  filter_out_expected[2793] <= 8'hfe;
  filter_out_expected[2794] <= 8'hfd;
  filter_out_expected[2795] <= 8'hf9;
  filter_out_expected[2796] <= 8'hf7;
  filter_out_expected[2797] <= 8'hf4;
  filter_out_expected[2798] <= 8'hef;
  filter_out_expected[2799] <= 8'hed;
  filter_out_expected[2800] <= 8'hee;
  filter_out_expected[2801] <= 8'hf2;
  filter_out_expected[2802] <= 8'hf8;
  filter_out_expected[2803] <= 8'hfe;
  filter_out_expected[2804] <= 8'hff;
  filter_out_expected[2805] <= 8'hfe;
  filter_out_expected[2806] <= 8'hfe;
  filter_out_expected[2807] <= 8'hff;
  filter_out_expected[2808] <= 8'h00;
  filter_out_expected[2809] <= 8'hfb;
  filter_out_expected[2810] <= 8'hf3;
  filter_out_expected[2811] <= 8'hf0;
  filter_out_expected[2812] <= 8'hf5;
  filter_out_expected[2813] <= 8'hfd;
  filter_out_expected[2814] <= 8'h03;
  filter_out_expected[2815] <= 8'h06;
  filter_out_expected[2816] <= 8'h06;
  filter_out_expected[2817] <= 8'h08;
  filter_out_expected[2818] <= 8'h0a;
  filter_out_expected[2819] <= 8'h0c;
  filter_out_expected[2820] <= 8'h0c;
  filter_out_expected[2821] <= 8'h07;
  filter_out_expected[2822] <= 8'hfe;
  filter_out_expected[2823] <= 8'hf8;
  filter_out_expected[2824] <= 8'hf6;
  filter_out_expected[2825] <= 8'hfb;
  filter_out_expected[2826] <= 8'h00;
  filter_out_expected[2827] <= 8'h04;
  filter_out_expected[2828] <= 8'h05;
  filter_out_expected[2829] <= 8'h06;
  filter_out_expected[2830] <= 8'h05;
  filter_out_expected[2831] <= 8'h03;
  filter_out_expected[2832] <= 8'h04;
  filter_out_expected[2833] <= 8'h04;
  filter_out_expected[2834] <= 8'h03;
  filter_out_expected[2835] <= 8'hfd;
  filter_out_expected[2836] <= 8'hf9;
  filter_out_expected[2837] <= 8'hfb;
  filter_out_expected[2838] <= 8'h04;
  filter_out_expected[2839] <= 8'h0a;
  filter_out_expected[2840] <= 8'h0a;
  filter_out_expected[2841] <= 8'h07;
  filter_out_expected[2842] <= 8'h04;
  filter_out_expected[2843] <= 8'h02;
  filter_out_expected[2844] <= 8'h01;
  filter_out_expected[2845] <= 8'h00;
  filter_out_expected[2846] <= 8'h03;
  filter_out_expected[2847] <= 8'h04;
  filter_out_expected[2848] <= 8'h01;
  filter_out_expected[2849] <= 8'hfe;
  filter_out_expected[2850] <= 8'hfc;
  filter_out_expected[2851] <= 8'hff;
  filter_out_expected[2852] <= 8'h01;
  filter_out_expected[2853] <= 8'hff;
  filter_out_expected[2854] <= 8'hfc;
  filter_out_expected[2855] <= 8'hff;
  filter_out_expected[2856] <= 8'h07;
  filter_out_expected[2857] <= 8'h11;
  filter_out_expected[2858] <= 8'h10;
  filter_out_expected[2859] <= 8'h08;
  filter_out_expected[2860] <= 8'h04;
  filter_out_expected[2861] <= 8'h03;
  filter_out_expected[2862] <= 8'h08;
  filter_out_expected[2863] <= 8'h08;
  filter_out_expected[2864] <= 8'h07;
  filter_out_expected[2865] <= 8'h07;
  filter_out_expected[2866] <= 8'h0a;
  filter_out_expected[2867] <= 8'h0a;
  filter_out_expected[2868] <= 8'h07;
  filter_out_expected[2869] <= 8'h02;
  filter_out_expected[2870] <= 8'hfd;
  filter_out_expected[2871] <= 8'hfa;
  filter_out_expected[2872] <= 8'hfb;
  filter_out_expected[2873] <= 8'hff;
  filter_out_expected[2874] <= 8'h02;
  filter_out_expected[2875] <= 8'h05;
  filter_out_expected[2876] <= 8'h02;
  filter_out_expected[2877] <= 8'h00;
  filter_out_expected[2878] <= 8'h05;
  filter_out_expected[2879] <= 8'h0a;
  filter_out_expected[2880] <= 8'h0f;
  filter_out_expected[2881] <= 8'h0e;
  filter_out_expected[2882] <= 8'h0a;
  filter_out_expected[2883] <= 8'h03;
  filter_out_expected[2884] <= 8'hfc;
  filter_out_expected[2885] <= 8'hf9;
  filter_out_expected[2886] <= 8'hfd;
  filter_out_expected[2887] <= 8'h03;
  filter_out_expected[2888] <= 8'h08;
  filter_out_expected[2889] <= 8'h09;
  filter_out_expected[2890] <= 8'h07;
  filter_out_expected[2891] <= 8'h03;
  filter_out_expected[2892] <= 8'h00;
  filter_out_expected[2893] <= 8'hfb;
  filter_out_expected[2894] <= 8'hf7;
  filter_out_expected[2895] <= 8'hf6;
  filter_out_expected[2896] <= 8'hf8;
  filter_out_expected[2897] <= 8'hfb;
  filter_out_expected[2898] <= 8'hfd;
  filter_out_expected[2899] <= 8'hfe;
  filter_out_expected[2900] <= 8'hfe;
  filter_out_expected[2901] <= 8'hfe;
  filter_out_expected[2902] <= 8'hfb;
  filter_out_expected[2903] <= 8'hf5;
  filter_out_expected[2904] <= 8'hf0;
  filter_out_expected[2905] <= 8'hf1;
  filter_out_expected[2906] <= 8'hf4;
  filter_out_expected[2907] <= 8'hf9;
  filter_out_expected[2908] <= 8'hf9;
  filter_out_expected[2909] <= 8'hf6;
  filter_out_expected[2910] <= 8'hf7;
  filter_out_expected[2911] <= 8'hfe;
  filter_out_expected[2912] <= 8'h02;
  filter_out_expected[2913] <= 8'h05;
  filter_out_expected[2914] <= 8'h04;
  filter_out_expected[2915] <= 8'h00;
  filter_out_expected[2916] <= 8'h01;
  filter_out_expected[2917] <= 8'h06;
  filter_out_expected[2918] <= 8'h09;
  filter_out_expected[2919] <= 8'h06;
  filter_out_expected[2920] <= 8'h01;
  filter_out_expected[2921] <= 8'hfd;
  filter_out_expected[2922] <= 8'hff;
  filter_out_expected[2923] <= 8'h03;
  filter_out_expected[2924] <= 8'h06;
  filter_out_expected[2925] <= 8'h03;
  filter_out_expected[2926] <= 8'hff;
  filter_out_expected[2927] <= 8'h01;
  filter_out_expected[2928] <= 8'h07;
  filter_out_expected[2929] <= 8'h0a;
  filter_out_expected[2930] <= 8'h0a;
  filter_out_expected[2931] <= 8'h05;
  filter_out_expected[2932] <= 8'h04;
  filter_out_expected[2933] <= 8'h02;
  filter_out_expected[2934] <= 8'h00;
  filter_out_expected[2935] <= 8'hfe;
  filter_out_expected[2936] <= 8'hfb;
  filter_out_expected[2937] <= 8'hfa;
  filter_out_expected[2938] <= 8'hfe;
  filter_out_expected[2939] <= 8'h02;
  filter_out_expected[2940] <= 8'h03;
  filter_out_expected[2941] <= 8'h03;
  filter_out_expected[2942] <= 8'hfe;
  filter_out_expected[2943] <= 8'hfa;
  filter_out_expected[2944] <= 8'hfb;
  filter_out_expected[2945] <= 8'hfc;
  filter_out_expected[2946] <= 8'hfe;
  filter_out_expected[2947] <= 8'h01;
  filter_out_expected[2948] <= 8'h02;
  filter_out_expected[2949] <= 8'h01;
  filter_out_expected[2950] <= 8'h02;
  filter_out_expected[2951] <= 8'h05;
  filter_out_expected[2952] <= 8'h0a;
  filter_out_expected[2953] <= 8'h0c;
  filter_out_expected[2954] <= 8'h07;
  filter_out_expected[2955] <= 8'h01;
  filter_out_expected[2956] <= 8'hfc;
  filter_out_expected[2957] <= 8'hfa;
  filter_out_expected[2958] <= 8'hfc;
  filter_out_expected[2959] <= 8'h02;
  filter_out_expected[2960] <= 8'h09;
  filter_out_expected[2961] <= 8'h10;
  filter_out_expected[2962] <= 8'h0f;
  filter_out_expected[2963] <= 8'h09;
  filter_out_expected[2964] <= 8'h03;
  filter_out_expected[2965] <= 8'h03;
  filter_out_expected[2966] <= 8'h06;
  filter_out_expected[2967] <= 8'h09;
  filter_out_expected[2968] <= 8'h08;
  filter_out_expected[2969] <= 8'h08;
  filter_out_expected[2970] <= 8'h08;
  filter_out_expected[2971] <= 8'h06;
  filter_out_expected[2972] <= 8'h04;
  filter_out_expected[2973] <= 8'hff;
  filter_out_expected[2974] <= 8'hfd;
  filter_out_expected[2975] <= 8'hfa;
  filter_out_expected[2976] <= 8'hf8;
  filter_out_expected[2977] <= 8'hf8;
  filter_out_expected[2978] <= 8'hfc;
  filter_out_expected[2979] <= 8'h00;
  filter_out_expected[2980] <= 8'h05;
  filter_out_expected[2981] <= 8'h06;
  filter_out_expected[2982] <= 8'h03;
  filter_out_expected[2983] <= 8'hff;
  filter_out_expected[2984] <= 8'hfb;
  filter_out_expected[2985] <= 8'hf9;
  filter_out_expected[2986] <= 8'hfb;
  filter_out_expected[2987] <= 8'hfe;
  filter_out_expected[2988] <= 8'h02;
  filter_out_expected[2989] <= 8'h07;
  filter_out_expected[2990] <= 8'h0b;
  filter_out_expected[2991] <= 8'h08;
  filter_out_expected[2992] <= 8'h05;
  filter_out_expected[2993] <= 8'h04;
  filter_out_expected[2994] <= 8'h06;
  filter_out_expected[2995] <= 8'h05;
  filter_out_expected[2996] <= 8'h01;
  filter_out_expected[2997] <= 8'hfa;
  filter_out_expected[2998] <= 8'hf8;
  filter_out_expected[2999] <= 8'hf9;
  filter_out_expected[3000] <= 8'hfa;
  filter_out_expected[3001] <= 8'hfb;
  filter_out_expected[3002] <= 8'hfe;
  filter_out_expected[3003] <= 8'h02;
  filter_out_expected[3004] <= 8'h04;
  filter_out_expected[3005] <= 8'h03;
  filter_out_expected[3006] <= 8'hff;
  filter_out_expected[3007] <= 8'hfd;
  filter_out_expected[3008] <= 8'hfe;
  filter_out_expected[3009] <= 8'h05;
  filter_out_expected[3010] <= 8'h07;
  filter_out_expected[3011] <= 8'h08;
  filter_out_expected[3012] <= 8'h05;
  filter_out_expected[3013] <= 8'h05;
  filter_out_expected[3014] <= 8'h03;
  filter_out_expected[3015] <= 8'h00;
  filter_out_expected[3016] <= 8'hfc;
  filter_out_expected[3017] <= 8'hfa;
  filter_out_expected[3018] <= 8'hfa;
  filter_out_expected[3019] <= 8'hfb;
  filter_out_expected[3020] <= 8'h00;
  filter_out_expected[3021] <= 8'h04;
  filter_out_expected[3022] <= 8'h0b;
  filter_out_expected[3023] <= 8'h0b;
  filter_out_expected[3024] <= 8'h07;
  filter_out_expected[3025] <= 8'h02;
  filter_out_expected[3026] <= 8'hfe;
  filter_out_expected[3027] <= 8'hfc;
  filter_out_expected[3028] <= 8'hfe;
  filter_out_expected[3029] <= 8'h01;
  filter_out_expected[3030] <= 8'h02;
  filter_out_expected[3031] <= 8'h03;
  filter_out_expected[3032] <= 8'h02;
  filter_out_expected[3033] <= 8'h05;
  filter_out_expected[3034] <= 8'h07;
  filter_out_expected[3035] <= 8'h05;
  filter_out_expected[3036] <= 8'h01;
  filter_out_expected[3037] <= 8'hfe;
  filter_out_expected[3038] <= 8'hfd;
  filter_out_expected[3039] <= 8'hfb;
  filter_out_expected[3040] <= 8'hfb;
  filter_out_expected[3041] <= 8'hfc;
  filter_out_expected[3042] <= 8'hfd;
  filter_out_expected[3043] <= 8'hfb;
  filter_out_expected[3044] <= 8'hf4;
  filter_out_expected[3045] <= 8'hf1;
  filter_out_expected[3046] <= 8'hf7;
  filter_out_expected[3047] <= 8'hff;
  filter_out_expected[3048] <= 8'h03;
  filter_out_expected[3049] <= 8'h00;
  filter_out_expected[3050] <= 8'hfe;
  filter_out_expected[3051] <= 8'hfd;
  filter_out_expected[3052] <= 8'hfd;
  filter_out_expected[3053] <= 8'hfd;
  filter_out_expected[3054] <= 8'hfd;
  filter_out_expected[3055] <= 8'hfc;
  filter_out_expected[3056] <= 8'hff;
  filter_out_expected[3057] <= 8'h03;
  filter_out_expected[3058] <= 8'h07;
  filter_out_expected[3059] <= 8'h08;
  filter_out_expected[3060] <= 8'h04;
  filter_out_expected[3061] <= 8'hfd;
  filter_out_expected[3062] <= 8'hf6;
  filter_out_expected[3063] <= 8'hf7;
  filter_out_expected[3064] <= 8'hfc;
  filter_out_expected[3065] <= 8'hff;
  filter_out_expected[3066] <= 8'h00;
  filter_out_expected[3067] <= 8'hfd;
  filter_out_expected[3068] <= 8'hfa;
  filter_out_expected[3069] <= 8'hfc;
  filter_out_expected[3070] <= 8'h00;
  filter_out_expected[3071] <= 8'h02;
  filter_out_expected[3072] <= 8'h04;
  filter_out_expected[3073] <= 8'h03;
  filter_out_expected[3074] <= 8'h00;
  filter_out_expected[3075] <= 8'hfb;
  filter_out_expected[3076] <= 8'hf6;
  filter_out_expected[3077] <= 8'hf5;
  filter_out_expected[3078] <= 8'hf6;
  filter_out_expected[3079] <= 8'hfb;
  filter_out_expected[3080] <= 8'h00;
  filter_out_expected[3081] <= 8'h08;
  filter_out_expected[3082] <= 8'h0c;
  filter_out_expected[3083] <= 8'h0b;
  filter_out_expected[3084] <= 8'h02;
  filter_out_expected[3085] <= 8'hfe;
  filter_out_expected[3086] <= 8'hff;
  filter_out_expected[3087] <= 8'h05;
  filter_out_expected[3088] <= 8'h09;
  filter_out_expected[3089] <= 8'h06;
  filter_out_expected[3090] <= 8'h01;
  filter_out_expected[3091] <= 8'hfd;
  filter_out_expected[3092] <= 8'hff;
  filter_out_expected[3093] <= 8'hff;
  filter_out_expected[3094] <= 8'hfe;
  filter_out_expected[3095] <= 8'hfa;
  filter_out_expected[3096] <= 8'hf9;
  filter_out_expected[3097] <= 8'hf8;
  filter_out_expected[3098] <= 8'hfa;
  filter_out_expected[3099] <= 8'hfc;
  filter_out_expected[3100] <= 8'h00;
  filter_out_expected[3101] <= 8'h02;
  filter_out_expected[3102] <= 8'h04;
  filter_out_expected[3103] <= 8'h02;
  filter_out_expected[3104] <= 8'h00;
  filter_out_expected[3105] <= 8'hff;
  filter_out_expected[3106] <= 8'h00;

  end // Input & Output data
//************************************


  parameter MAX_TIMEOUT = 3; //uint32
  parameter MAX_ERROR_COUNT = 3107; //uint32


 // Signals
  reg  clk; // boolean
  reg  clk_enable; // boolean
  reg  syn_rst; // boolean
  reg  signed [7:0] filter_in; // sfix8_En7
  wire signed [7:0] filter_out; // sfix8_En7

  reg  tb_enb; // boolean
  wire srcDone; // boolean
  wire snkDone; // boolean
  wire testFailure; // boolean
  reg  tbenb_dly; // boolean
  reg  rdEnb; // boolean
  wire filter_in_data_log_rdenb; // boolean
  reg  [11:0] filter_in_data_log_addr; // ufix12
  reg  filter_in_data_log_done; // boolean
  reg  filter_out_testFailure; // boolean
  integer filter_out_timeout; // uint32
  integer filter_out_errCnt; // uint32
  wire delayLine_out; // boolean
  wire expected_ce_out; // boolean
  reg  int_delay_pipe [0:1] ; // boolean
  wire filter_out_rdenb; // boolean
  reg  [11:0] filter_out_addr; // ufix12
  reg  filter_out_done; // boolean
  wire signed [7:0] filter_out_ref; // sfix8_En7
  reg  check1_Done; // boolean

 // Module Instances
  fir_da u_fir_da
    (
    .clk(clk),
    .clk_enable(clk_enable),
    .syn_rst(syn_rst),
    .filter_in(filter_in),
    .filter_out(filter_out)
    );


 // Block Statements
  // -------------------------------------------------------------
  // Driving the test bench enable
  // -------------------------------------------------------------

  always @(syn_rst, snkDone)
  begin
    if (syn_rst == 1'b1)
      tb_enb <= 1'b0;
    else if (snkDone == 1'b0 )
      tb_enb <= 1'b1;
    else begin
    # (clk_period * 2);
      tb_enb <= 1'b0;
    end
  end

  always @(posedge clk or posedge syn_rst) // completed_msg
  begin
    if (syn_rst) begin 
       // Nothing to reset.
    end 
    else begin 
      if (snkDone == 1) begin
        if (testFailure == 0)
              $display("**************TEST COMPLETED (PASSED)**************");
        else
              $display("**************TEST COMPLETED (FAILED)**************");
      end
    end
  end // completed_msg;

  // -------------------------------------------------------------
  // System Clock (fast clock) and reset
  // -------------------------------------------------------------

  always  // clock generation
  begin // clk_gen
    clk <= 1'b1;
    # clk_high;
    clk <= 1'b0;
    # clk_low;
    if (snkDone == 1) begin
      clk <= 1'b1;
      # clk_high;
      clk <= 1'b0;
      # clk_low;
      $stop;
    end
  end  // clk_gen

  initial  // reset block
  begin // syn_rst_gen
    syn_rst <= 1'b1;
    # (clk_period * 2);
    @ (posedge clk);
    # (clk_hold);
    syn_rst <= 1'b0;
  end  // syn_rst_gen

  // -------------------------------------------------------------
  // Testbench clock enable
  // -------------------------------------------------------------

  always @ ( posedge clk)
    begin: tb_enb_delay
      if (syn_rst == 1'b1) begin
        tbenb_dly <= 1'b0;
      end
      else begin
        if (tb_enb == 1'b1) begin
          tbenb_dly <= tb_enb;
        end
      end
    end // tb_enb_delay

  always @(snkDone, tbenb_dly)
  begin
    if (snkDone == 0)
      rdEnb <= tbenb_dly;
    else
      rdEnb <= 0;
  end

  // -------------------------------------------------------------
  // Read the data and transmit it to the DUT
  // -------------------------------------------------------------

  always @(posedge clk or posedge syn_rst)
  begin
    filter_in_data_log_task(clk,syn_rst,
                            filter_in_data_log_rdenb,filter_in_data_log_addr,
                            filter_in_data_log_done);
  end

  assign filter_in_data_log_rdenb = rdEnb;

  always @ (filter_in_data_log_rdenb, filter_in_data_log_addr)
  begin // stimuli_filter_in_data_log_filter_in
    if (filter_in_data_log_rdenb == 1) begin
      filter_in <= # clk_hold filter_in_data_log_force[filter_in_data_log_addr];
    end
  end // stimuli_filter_in_data_log_filter_in

  // -------------------------------------------------------------
  // Create done signal for Input data
  // -------------------------------------------------------------

  assign srcDone = filter_in_data_log_done;


  always @( posedge clk)
    begin: ceout_delayLine
      if (syn_rst == 1'b1) begin
        int_delay_pipe[0] <= 1'b0;
        int_delay_pipe[1] <= 1'b0;
      end
      else begin
        if (clk_enable == 1'b1) begin
        int_delay_pipe[0] <= rdEnb;
        int_delay_pipe[1] <= int_delay_pipe[0];
        end
      end
    end // ceout_delayLine

  assign delayLine_out = int_delay_pipe[1];

  assign expected_ce_out =  delayLine_out & clk_enable;

  // -------------------------------------------------------------
  //  Checker: Checking the data received from the DUT.
  // -------------------------------------------------------------

  always @(posedge clk or posedge syn_rst)
  begin
    filter_out_task(clk,syn_rst,
                    filter_out_rdenb,filter_out_addr,
                    filter_out_done);
  end

  assign filter_out_rdenb = expected_ce_out;

  assign filter_out_ref = filter_out_expected[filter_out_addr];


  always @ (posedge clk or posedge syn_rst) // checker_filter_out
  begin
    if (syn_rst == 1) begin
      filter_out_timeout <= 0;
      filter_out_testFailure <= 0;
      filter_out_errCnt <= 0;
    end 
    else begin 
      if (filter_out_rdenb == 1 ) begin 
        filter_out_timeout <= 0;
        if (((abs(filter_out - filter_out_expected[filter_out_addr]) > 15) !== 0 )) begin
           filter_out_errCnt <= filter_out_errCnt + 1;
           filter_out_testFailure <= 1;
                   $display("ERROR  in filter_out at time %t : Expected '%h' Actual '%h'", 
                        $time, filter_out_expected[filter_out_addr], filter_out);
           if (filter_out_errCnt >= MAX_ERROR_COUNT) 
             $display("Warning: Number of errors for filter_out have exceeded the maximum error limit");
        end

      end
      else if (filter_out_timeout > MAX_TIMEOUT && filter_out_rdenb == 1 ) begin 
        filter_out_errCnt <= filter_out_errCnt + 1;
        filter_out_testFailure <= 1;
        $display ("Error: Timeout - Data was not received for filter_out.");
        $stop;
      end
      else if (filter_out_rdenb == 1) begin
        filter_out_timeout <= filter_out_timeout + 1 ;
      end
    end
  end // checker_filter_out

  always @ (posedge clk or posedge syn_rst) // checkDone_1
  begin
    if (syn_rst == 1)
      check1_Done <= 0;
    else if ((check1_Done == 0) && (filter_out_done == 1) && (filter_out_rdenb == 1))
      check1_Done <= 1;
  end

  // -------------------------------------------------------------
  // Create done and test failure signal for output data
  // -------------------------------------------------------------

  assign snkDone = check1_Done;

  assign testFailure = filter_out_testFailure;

  // -------------------------------------------------------------
  // Global clock enable
  // -------------------------------------------------------------
  always @(snkDone, tbenb_dly)
  begin
    if (snkDone == 0)
      # clk_hold clk_enable <= tbenb_dly;
    else
      # clk_hold clk_enable <= 0;
  end

 // Assignment Statements



endmodule // filter_tb
