
--------------------------------------------
-- Architecture
--------------------------------------------
architecture rtl of wiener_coeff is

  type ROM_STORAGE_T is array (0 to 2**(WIENER_ADDR_WIDTH_CT)-1) of
                     std_logic_vector((4*WIENER_COEFF_WIDTH_CT)-1 downto 0);
                     
  -----------------------------------------------------------------------------
  -- array only requires 0 to 287 locations, but CVE fails by testing addresses
  -- greater than that (which is prevented in reality by the logic)
  -- Therefore, increased the size of the array and used an others clause.
  -----------------------------------------------------------------------------
  constant WIENER_COEFF_CT : ROM_STORAGE_T := (
              "1111111110111101001000001101010111101011",
              "1111111100111111000000000000110000011000",
              "0000000101111111010000000001000000001100",
              "1111011001001010100001011001010000110101",
              "1111111100000010011100000100001111000100",
              "1111110100000001011100000000011111100011",
              "0010100000010000011000101010001111010010",
              "0000011100111111011011110011010000000110",
              "0000000100000000000111111011010000001001",
              "0100000110001010000011110110011111111110",
              "1111110110111100100000000001100010100101",
              "0000001100111110001100000010010000100010",
              "0010100101000000011011110001000000011000",
              "1111001110000000111100101000000011110010",
              "1111111100111111110000000111001111110110",
              "0000000110111100110100000100000000000011",
              "0000001111001010010100111100110010100000",
              "1111110000000010011111111101101111001000",
              "1111111101111100101000000110011111111111",
              "1111111101001010001100111111110010100011",
              "0000000000111111111100000110011111001010",
              "1111111110111100110100000101100000000000",
              "1111111111001010100100111111010010011111",
              "1111111110000000000000001000001110111110",
              "0000000101111100111000000100000000000011",
              "0000001110001010011100111100110010011111",
              "1111110010000010000000000000001111000001",
              "1111111110111100101100000101100000000000",
              "1111101001001010010000111111110010100010",
              "1111110001000011000011110100100000000000",
              "0000000101111100111000000100000000000011",
              "0000000000001010111000111101000010011101",
              "1111110001000010010011111101101111010001",
              "1111100011111100011000001010001111111001",
              "0001110001000000000001010110000010101001",
              "1111110010000011000111110101101111001011",
              "1111001011111101011000001100011111110010",
              "0010101001010101100000000000000001110001",
              "1111111001000010100011110001101111100011",
              "1111010001111111011000001001001111110001",
              "0010011101001111010000101011100000000000",
              "0000000011000001000011110011100000000101",
              "0000000000111101001000001100001111110001",
              "0010100010001111111100101001001111101001",
              "0000000000000001011011110010111111111110",
              "1111000001000000000000001000001111110010",
              "0010011111001111001100101001110000001110",
              "0000000011000001000011110011100000000101",
              "1110111110000010000000000000001111111110",
              "0010011111001111110100101010011111111111",
              "0000000000000001011011110011011111111110",
              "1111001010000001100111111111110000000000",
              "0010100011001111111100101000111111111101",
              "1111111111000001100111110010101111111101",
              "1111001000111111011000001001111111110000",
              "0010100000001111001100101001010000001111",
              "0000000011000001000011110011010000000110",
              "1111110110000001110011111111001111111100",
              "0011110010001010000000000011111111001110",
              "0000011000111100010000000001100010100101",
              "0000100010000000100111111000110000001100",
              "0010100101000000011011110010001111110110",
              "1111111110111101100100101000000100000110",
              "0000001001111110110100000000010000000100",
              "0000000110111100110111111101100000011100",
              "1111010010001010100001000001100010100000",
              "1111100011000000000100000101111111110100",
              "1111000100000001000000001001111111111100",
              "0000110101010110010100101010001111011001",
              "0000001100000000010011111101000000000101",
              "0000011000000000001111111100001111111100",
              "0111101011000011010111110100101111111110",
              "1111011111111101001100010110100111011000",
              "1111110000000000011100000110100000001100",
              "1111110111000001000000000001101111110001",
              "0000011100001011100101000100110001011010",
              "0000100011000000101011110101011111001000",
              "0000010000111110110011111011000000001110",
              "0010010110001110100000101110011111010011",
              "0000000011111101111111110111110000100011",
              "0000000110111110110000000001110000011000",
              "0011001110001001011000000111001111011111",
              "1111010110111110010100001101100010011110",
              "1111110001000000111000000110001111111001",
              "0010011110000010001111110010000000001100",
              "1111100000000011001000100111000011010000",
              "1111110000000010001100000000111111010110",
              "0000110110111101111111110101010000011010",
              "0000110010001001010100110001010010011100",
              "0000000111000000101011110111111111100101",
              "0000110100111110000011110110000000011001",
              "0000110100001001100100110001100010011001",
              "0000000000000001100111110110001111100000",
              "0000110111111101111011110101000000011011",
              "0000110000001001001100110001010010011101",
              "0000001010000000000011111001111111100110",
              "0000110100111101111011110110000000011001",
              "0000101110001001100100110010010010011011",
              "0000001100111111010000000000001111010100",
              "0000110111111101110111110101000000011011",
              "0000100100001001000000110001110010100000",
              "0000001010000000011111110100100000000000",
              "0000110000111101111111110110110000011000",
              "0000000000001010111100110011010010010111",
              "0000001001000000000111111001011111111111",
              "0000101010111100111111110110100000011101",
              "0001111100000000000001000010110010110100",
              "0000010011111111011011110011111111111111",
              "1111111111111100111111111101100000010011",
              "0010110100010000101100000000000001111100",
              "0000011101111101101011110011110000101010",
              "1111111111111110010100000000010000001001",
              "0010010111001100110100101011110000000000",
              "0000011000111101101111110111110000110000",
              "0000000000111101001000000001110000001010",
              "0010100000001100011100100100000000100100",
              "0000011011111101010011110111010000110111",
              "1111010100000000000011111101000000001100",
              "0010011011001100100100100110010000101110",
              "0000011001111101100011110111100000110100",
              "1111100110111110011100000000000000001010",
              "0010011101001100010100100100110000110000",
              "0000011011111101010011110111100000110111",
              "1111100000111101100000000110010000000000",
              "0010011001001100011000100110010000110100",
              "0000011001111101100011111000000000110100",
              "1111100101111101111100000010100000000111",
              "0010011100001100010100100101010000110010",
              "0000011010111101010111110111110000110110",          
              "1111010110000000001100001000111111110000",
              "0011010000001001110000001100101111100000",
              "0000001100111100100000001000110010011110",
              "1111111001000001100000000011101111110001",
              "0010011110000011011011111001011111010110",
              "1111011111000001110000100101100011001110",
              "0000011000000000011111111011000000000110",
              "0000100011111101111111110111110000000011",
              "1111010011001011100100111010000010010110",
              "0000001110111110110011111011000000010000",
              "1111001000111101010100000010100000100011",
              "0001011010010001001100101110010000011100",
              "1111110001000000011000000100001111110111",
              "0000001100000001101000000001111111110000",
              "0111011000000101101011110100111111011111",
              "1111011000000001010100101000100110010001",
              "0000010101000000010011111010001111010010",
              "1111110110111111100000000010000000010110",
              "0001001111001000010000101001110010100010",
              "1111100111111110001011111100100000011001",
              "1111111000000001001000000011101111111010",
              "0010001011001010010000100001000000010101",
              "1111100000111111000100000111000001010110",
              "0000001000000000111011111111001111100110",
              "0010010110001000101100010011111111011000",
              "1111110111000001111000010011100001111100",
              "0000010110111111101011111001101111100100",
              "0001111100000101011000000110011111010010",
              "0000100010000101000100011101100010000111",
              "0000010101111110011111111000001111110111",
              "0001001110000001110011111100101111101000",
              "0001010001000111100000100001100001110110",
              "0000000100111110001011111100010000011110",
              "0001001111000001110011111100101111101000",
              "0001001111000111011100100001100001110111",
              "0000000000111110100011111100100000011100",
              "0001001111000001101111111100011111101001",
              "0001001111000111100100100010000001111000",
              "1111110110000000000011111001100000010111",
              "0001001111000001110011111100101111101000",
              "0001001101000111011100100001100001110111",
              "0000000011111101110000000000000000011000",
              "0001001100000001101011111100101111101010",
              "0001011011000111111000100010000001110101",
              "0000000001111110100011111111010000000000",
              "0001001101000001010111111011011111101101",
              "0000000000001001000100100101110001111101",
              "1111111010111110011100000001000000111000",
              "0001011000000001011111111010011111101001",
              "0001110110000000000000101010110010010000",
              "1111111100111101111011111110100000110111",
              "0000110111111111101011110111101111111100",
              "0010010000001010101100000000000001110110",
              "1111101001111110100100000101110001011000",
              "0000111000000000010011111001111111111010",
              "0001111101001001011100100100010000000000",
              "1111101101111110110100000101010001001101",
              "0000000000111111110111111010000000000001",
              "0001110101001000100000011111100001011011",
              "1111101010111111001000000110100001001100",
              "0000011000000000000011110111000000000011",
              "0001110111001000011000011101110001001101",
              "1111101000111111001000000111000001001111",
              "0000010111111110011000000000001111110110",
              "0001111000001000100000011110010001001111",
              "1111101001111111000100000110110001001111",
              "0000011100111111001011111010000000000000",
              "0001110111001000011000011101110001001111",
              "1111101000111111001000000111000001001111",
              "0000011110111111000111111000100000000100",
              "0001110110001000011000011110000001010001",
              "1111101000111111001000000111000001001110",
              "1111110111111110000011111001110000010101",
              "0010000111000111011000010100010000100010",
              "1111010010000001100100010101100001111100",
              "1111100100111110011011111110100000010110",
              "0001111100000100111000000111101111110111",
              "1111011000000100111100100010110010010110",
              "1111100110111111110000000011100000001000",
              "0001010110000001110011111100011111100000",
              "0000010101001000010000101001000010001011",
              "1111111010000000111000000100101111111000",
              "0000011001111111001011111000101111100111",
              "0010100010001010011100100001000001001111",
              "0000010110000000100011111110001111110110",
              "1111010010111110100000000001000000010101",
              "0110010001001010001000000101011111011000",
              "0000010010000101011000101110000100111101",
              "1111100101111101101011110110011111101010",
              "0000001111000001000100000010001111110111",
              "0001000101000110100100100100000010111000",
              "1111110000111111101100000011010000100110",
              "0000010001111111111011111100011111101100",
              "0001100001000110110000011010010001010110",
              "0000000011000001101000001101010001001110",
              "0000001000111111000111111010111111110010",
              "0001101010000110000100010001010000010010",
              "0000011011000011011100010100000001100011",
              "1111110111111110110011111100100000000011",
              "0001100011000100111000001001101111101010",
              "0000110110000100111000011000000001101000",
              "1111100101111111000000000000110000011011",
              "0001010000000011010100000011011111011001",
              "0001001110000101111000011001000001100000",
              "1111011010111111101100000110100000110111",
              "0001010010000011001100000010011111010110",
              "0001010010000110010100011011000001100101",
              "0000000000111101011000000010010000110011",
              "0001010001000011010100000011011111011001",
              "0001001101000101110100011001000001100000",
              "1111010111000000000000000110010000110110",
              "0001001111000011001100000011001111011010",
              "0001010011000110000100011001100001100000",
              "1111011111000000000100000000000000111101",
              "0001010001000011001100000010101111011000",
              "0001011011000110100000011010110001100100",
              "1111011100000000010000001010000000000000",
              "0001010110000011010100000010101111010100",
              "0000000000000111000000011100110001101010",
              "1111010101000000001000001010010001001010",
              "0001011101000011101100000011001111010000",
              "0001100100000000000000011110010001110010",
              "1111010001111111110100001001100001001001",
              "0001001001000010011011111111011111010001",
              "0001110010000111100100000000000001100100",
              "1111010000000000110000001110110001011101",
              "0001001010000010100100000000101111010101",
              "0001101010000111001100011100000000000000",
              "1111010100000000101000001101010001010110",
              "0000000000000010100000000001001111011100",
              "0001100100000110101100011010000001011011",
              "1111011000000000101000001100110001010001",
              "0000111101000000000000000000011111011111",
              "0001100000000110011000011000010001010011",
              "1111011010000000110000001100110001001111",
              "0000110110000001100100000000001111010111",
              "0001100000000110010000010111010001001101",
              "1111011001000000110100001101010001010001",
              "0000110011000000100111110101100000000000",
              "0001100101000110110000011001010001010010",
              "1111010110000000100100001100110001010010",
              "0000110111000001101011111110111111011010",
              "0001100000000110010000010111100001001110",
              "1111011001000000110100001101010001010000",
              "0000011011000000001111111100001111100101",
              "0001101000000110000000010011100000110110",
              "1111101010000010011000010011100001100011",
              "0000000011111111001011111011001111110111",
              "0001100011000101000000001101110000011011",
              "0000010010000100010100011000010001101010",
              "1111110010111110101111111100010000001000",
              "0001001110000011010100000110100000000011",
              "0001010110000110100100011011000001100001",
              "1111101100111111000111111111100000010001",
              "0000100110000000110111111110111111110000",
              "0010111000001001000000011010010001000101",
              "1111110111000000100000000100010000001111",
              "1111101010111101100111110110101111100101",
              "0100111101001011100000010101100000010010",
    others => "0100111101001011100000010101100000010010"
             );


begin

  --------------------------------------------
  -- Output the coefficient corresponding to the input address.
  --------------------------------------------
  registers_p: process (clk, reset_n)
    variable chanwien_a_int_v : 
                 integer range 0 to 2**(WIENER_ADDR_WIDTH_CT)-1;
  begin
    if reset_n = '0' then               -- asynchronous reset (active low)
      chanwien_do_o       <= (others => '0');
    elsif clk'event and clk = '1' then  -- rising clock edge
      if module_enable_i = '1' then
        chanwien_a_int_v := conv_integer(chanwien_a_i);
        if chanwien_cs_ni = '0' then
          chanwien_do_o <= WIENER_COEFF_CT(chanwien_a_int_v);
        end if;
      end if;
    end if;
  end process registers_p;

end rtl;
