

--------------------------------------------
-- Architecture
--------------------------------------------
architecture rtl of sine_table_rom is

  constant MAX_ADDR_CT : integer := 1024;

  type ROM_MEM_T is array (0 to MAX_ADDR_CT - 1) of integer ;
  
  signal sin_table : ROM_MEM_T ; -- sine table
  signal addr_tmp  : integer range MAX_ADDR_CT-1 downto 0 ; -- address
  signal sin_tmp   : std_logic_vector(9 downto 0); -- sine

begin

  -- sine table definition :
  sin_table(0) <= 0;
  sin_table(1) <= 2;
  sin_table(2) <= 3;
  sin_table(3) <= 5;
  sin_table(4) <= 6;
  sin_table(5) <= 8;
  sin_table(6) <= 9;
  sin_table(7) <= 11;
  sin_table(8) <= 13;
  sin_table(9) <= 14;
  sin_table(10) <= 16;
  sin_table(11) <= 17;
  sin_table(12) <= 19;
  sin_table(13) <= 20;
  sin_table(14) <= 22;
  sin_table(15) <= 24;
  sin_table(16) <= 25;
  sin_table(17) <= 27;
  sin_table(18) <= 28;
  sin_table(19) <= 30;
  sin_table(20) <= 31;
  sin_table(21) <= 33;
  sin_table(22) <= 35;
  sin_table(23) <= 36;
  sin_table(24) <= 38;
  sin_table(25) <= 39;
  sin_table(26) <= 41;
  sin_table(27) <= 42;
  sin_table(28) <= 44;
  sin_table(29) <= 45;
  sin_table(30) <= 47;
  sin_table(31) <= 49;
  sin_table(32) <= 50;
  sin_table(33) <= 52;
  sin_table(34) <= 53;
  sin_table(35) <= 55;
  sin_table(36) <= 56;
  sin_table(37) <= 58;
  sin_table(38) <= 60;
  sin_table(39) <= 61;
  sin_table(40) <= 63;
  sin_table(41) <= 64;
  sin_table(42) <= 66;
  sin_table(43) <= 67;
  sin_table(44) <= 69;
  sin_table(45) <= 71;
  sin_table(46) <= 72;
  sin_table(47) <= 74;
  sin_table(48) <= 75;
  sin_table(49) <= 77;
  sin_table(50) <= 78;
  sin_table(51) <= 80;
  sin_table(52) <= 82;
  sin_table(53) <= 83;
  sin_table(54) <= 85;
  sin_table(55) <= 86;
  sin_table(56) <= 88;
  sin_table(57) <= 89;
  sin_table(58) <= 91;
  sin_table(59) <= 92;
  sin_table(60) <= 94;
  sin_table(61) <= 96;
  sin_table(62) <= 97;
  sin_table(63) <= 99;
  sin_table(64) <= 100;
  sin_table(65) <= 102;
  sin_table(66) <= 103;
  sin_table(67) <= 105;
  sin_table(68) <= 107;
  sin_table(69) <= 108;
  sin_table(70) <= 110;
  sin_table(71) <= 111;
  sin_table(72) <= 113;
  sin_table(73) <= 114;
  sin_table(74) <= 116;
  sin_table(75) <= 117;
  sin_table(76) <= 119;
  sin_table(77) <= 121;
  sin_table(78) <= 122;
  sin_table(79) <= 124;
  sin_table(80) <= 125;
  sin_table(81) <= 127;
  sin_table(82) <= 128;
  sin_table(83) <= 130;
  sin_table(84) <= 131;
  sin_table(85) <= 133;
  sin_table(86) <= 135;
  sin_table(87) <= 136;
  sin_table(88) <= 138;
  sin_table(89) <= 139;
  sin_table(90) <= 141;
  sin_table(91) <= 142;
  sin_table(92) <= 144;
  sin_table(93) <= 145;
  sin_table(94) <= 147;
  sin_table(95) <= 149;
  sin_table(96) <= 150;
  sin_table(97) <= 152;
  sin_table(98) <= 153;
  sin_table(99) <= 155;
  sin_table(100) <= 156;
  sin_table(101) <= 158;
  sin_table(102) <= 159;
  sin_table(103) <= 161;
  sin_table(104) <= 163;
  sin_table(105) <= 164;
  sin_table(106) <= 166;
  sin_table(107) <= 167;
  sin_table(108) <= 169;
  sin_table(109) <= 170;
  sin_table(110) <= 172;
  sin_table(111) <= 173;
  sin_table(112) <= 175;
  sin_table(113) <= 176;
  sin_table(114) <= 178;
  sin_table(115) <= 180;
  sin_table(116) <= 181;
  sin_table(117) <= 183;
  sin_table(118) <= 184;
  sin_table(119) <= 186;
  sin_table(120) <= 187;
  sin_table(121) <= 189;
  sin_table(122) <= 190;
  sin_table(123) <= 192;
  sin_table(124) <= 193;
  sin_table(125) <= 195;
  sin_table(126) <= 196;
  sin_table(127) <= 198;
  sin_table(128) <= 200;
  sin_table(129) <= 201;
  sin_table(130) <= 203;
  sin_table(131) <= 204;
  sin_table(132) <= 206;
  sin_table(133) <= 207;
  sin_table(134) <= 209;
  sin_table(135) <= 210;
  sin_table(136) <= 212;
  sin_table(137) <= 213;
  sin_table(138) <= 215;
  sin_table(139) <= 216;
  sin_table(140) <= 218;
  sin_table(141) <= 220;
  sin_table(142) <= 221;
  sin_table(143) <= 223;
  sin_table(144) <= 224;
  sin_table(145) <= 226;
  sin_table(146) <= 227;
  sin_table(147) <= 229;
  sin_table(148) <= 230;
  sin_table(149) <= 232;
  sin_table(150) <= 233;
  sin_table(151) <= 235;
  sin_table(152) <= 236;
  sin_table(153) <= 238;
  sin_table(154) <= 239;
  sin_table(155) <= 241;
  sin_table(156) <= 242;
  sin_table(157) <= 244;
  sin_table(158) <= 246;
  sin_table(159) <= 247;
  sin_table(160) <= 249;
  sin_table(161) <= 250;
  sin_table(162) <= 252;
  sin_table(163) <= 253;
  sin_table(164) <= 255;
  sin_table(165) <= 256;
  sin_table(166) <= 258;
  sin_table(167) <= 259;
  sin_table(168) <= 261;
  sin_table(169) <= 262;
  sin_table(170) <= 264;
  sin_table(171) <= 265;
  sin_table(172) <= 267;
  sin_table(173) <= 268;
  sin_table(174) <= 270;
  sin_table(175) <= 271;
  sin_table(176) <= 273;
  sin_table(177) <= 274;
  sin_table(178) <= 276;
  sin_table(179) <= 277;
  sin_table(180) <= 279;
  sin_table(181) <= 280;
  sin_table(182) <= 282;
  sin_table(183) <= 283;
  sin_table(184) <= 285;
  sin_table(185) <= 286;
  sin_table(186) <= 288;
  sin_table(187) <= 289;
  sin_table(188) <= 291;
  sin_table(189) <= 292;
  sin_table(190) <= 294;
  sin_table(191) <= 295;
  sin_table(192) <= 297;
  sin_table(193) <= 298;
  sin_table(194) <= 300;
  sin_table(195) <= 301;
  sin_table(196) <= 303;
  sin_table(197) <= 304;
  sin_table(198) <= 306;
  sin_table(199) <= 307;
  sin_table(200) <= 309;
  sin_table(201) <= 310;
  sin_table(202) <= 312;
  sin_table(203) <= 313;
  sin_table(204) <= 315;
  sin_table(205) <= 316;
  sin_table(206) <= 318;
  sin_table(207) <= 319;
  sin_table(208) <= 321;
  sin_table(209) <= 322;
  sin_table(210) <= 324;
  sin_table(211) <= 325;
  sin_table(212) <= 327;
  sin_table(213) <= 328;
  sin_table(214) <= 330;
  sin_table(215) <= 331;
  sin_table(216) <= 333;
  sin_table(217) <= 334;
  sin_table(218) <= 336;
  sin_table(219) <= 337;
  sin_table(220) <= 339;
  sin_table(221) <= 340;
  sin_table(222) <= 342;
  sin_table(223) <= 343;
  sin_table(224) <= 345;
  sin_table(225) <= 346;
  sin_table(226) <= 348;
  sin_table(227) <= 349;
  sin_table(228) <= 351;
  sin_table(229) <= 352;
  sin_table(230) <= 353;
  sin_table(231) <= 355;
  sin_table(232) <= 356;
  sin_table(233) <= 358;
  sin_table(234) <= 359;
  sin_table(235) <= 361;
  sin_table(236) <= 362;
  sin_table(237) <= 364;
  sin_table(238) <= 365;
  sin_table(239) <= 367;
  sin_table(240) <= 368;
  sin_table(241) <= 370;
  sin_table(242) <= 371;
  sin_table(243) <= 373;
  sin_table(244) <= 374;
  sin_table(245) <= 375;
  sin_table(246) <= 377;
  sin_table(247) <= 378;
  sin_table(248) <= 380;
  sin_table(249) <= 381;
  sin_table(250) <= 383;
  sin_table(251) <= 384;
  sin_table(252) <= 386;
  sin_table(253) <= 387;
  sin_table(254) <= 389;
  sin_table(255) <= 390;
  sin_table(256) <= 391;
  sin_table(257) <= 393;
  sin_table(258) <= 394;
  sin_table(259) <= 396;
  sin_table(260) <= 397;
  sin_table(261) <= 399;
  sin_table(262) <= 400;
  sin_table(263) <= 402;
  sin_table(264) <= 403;
  sin_table(265) <= 404;
  sin_table(266) <= 406;
  sin_table(267) <= 407;
  sin_table(268) <= 409;
  sin_table(269) <= 410;
  sin_table(270) <= 412;
  sin_table(271) <= 413;
  sin_table(272) <= 415;
  sin_table(273) <= 416;
  sin_table(274) <= 417;
  sin_table(275) <= 419;
  sin_table(276) <= 420;
  sin_table(277) <= 422;
  sin_table(278) <= 423;
  sin_table(279) <= 425;
  sin_table(280) <= 426;
  sin_table(281) <= 427;
  sin_table(282) <= 429;
  sin_table(283) <= 430;
  sin_table(284) <= 432;
  sin_table(285) <= 433;
  sin_table(286) <= 435;
  sin_table(287) <= 436;
  sin_table(288) <= 437;
  sin_table(289) <= 439;
  sin_table(290) <= 440;
  sin_table(291) <= 442;
  sin_table(292) <= 443;
  sin_table(293) <= 444;
  sin_table(294) <= 446;
  sin_table(295) <= 447;
  sin_table(296) <= 449;
  sin_table(297) <= 450;
  sin_table(298) <= 452;
  sin_table(299) <= 453;
  sin_table(300) <= 454;
  sin_table(301) <= 456;
  sin_table(302) <= 457;
  sin_table(303) <= 459;
  sin_table(304) <= 460;
  sin_table(305) <= 461;
  sin_table(306) <= 463;
  sin_table(307) <= 464;
  sin_table(308) <= 466;
  sin_table(309) <= 467;
  sin_table(310) <= 468;
  sin_table(311) <= 470;
  sin_table(312) <= 471;
  sin_table(313) <= 473;
  sin_table(314) <= 474;
  sin_table(315) <= 475;
  sin_table(316) <= 477;
  sin_table(317) <= 478;
  sin_table(318) <= 479;
  sin_table(319) <= 481;
  sin_table(320) <= 482;
  sin_table(321) <= 484;
  sin_table(322) <= 485;
  sin_table(323) <= 486;
  sin_table(324) <= 488;
  sin_table(325) <= 489;
  sin_table(326) <= 491;
  sin_table(327) <= 492;
  sin_table(328) <= 493;
  sin_table(329) <= 495;
  sin_table(330) <= 496;
  sin_table(331) <= 497;
  sin_table(332) <= 499;
  sin_table(333) <= 500;
  sin_table(334) <= 502;
  sin_table(335) <= 503;
  sin_table(336) <= 504;
  sin_table(337) <= 506;
  sin_table(338) <= 507;
  sin_table(339) <= 508;
  sin_table(340) <= 510;
  sin_table(341) <= 511;
  sin_table(342) <= 512;
  sin_table(343) <= 514;
  sin_table(344) <= 515;
  sin_table(345) <= 516;
  sin_table(346) <= 518;
  sin_table(347) <= 519;
  sin_table(348) <= 521;
  sin_table(349) <= 522;
  sin_table(350) <= 523;
  sin_table(351) <= 525;
  sin_table(352) <= 526;
  sin_table(353) <= 527;
  sin_table(354) <= 529;
  sin_table(355) <= 530;
  sin_table(356) <= 531;
  sin_table(357) <= 533;
  sin_table(358) <= 534;
  sin_table(359) <= 535;
  sin_table(360) <= 537;
  sin_table(361) <= 538;
  sin_table(362) <= 539;
  sin_table(363) <= 541;
  sin_table(364) <= 542;
  sin_table(365) <= 543;
  sin_table(366) <= 545;
  sin_table(367) <= 546;
  sin_table(368) <= 547;
  sin_table(369) <= 549;
  sin_table(370) <= 550;
  sin_table(371) <= 551;
  sin_table(372) <= 553;
  sin_table(373) <= 554;
  sin_table(374) <= 555;
  sin_table(375) <= 557;
  sin_table(376) <= 558;
  sin_table(377) <= 559;
  sin_table(378) <= 560;
  sin_table(379) <= 562;
  sin_table(380) <= 563;
  sin_table(381) <= 564;
  sin_table(382) <= 566;
  sin_table(383) <= 567;
  sin_table(384) <= 568;
  sin_table(385) <= 570;
  sin_table(386) <= 571;
  sin_table(387) <= 572;
  sin_table(388) <= 574;
  sin_table(389) <= 575;
  sin_table(390) <= 576;
  sin_table(391) <= 577;
  sin_table(392) <= 579;
  sin_table(393) <= 580;
  sin_table(394) <= 581;
  sin_table(395) <= 583;
  sin_table(396) <= 584;
  sin_table(397) <= 585;
  sin_table(398) <= 586;
  sin_table(399) <= 588;
  sin_table(400) <= 589;
  sin_table(401) <= 590;
  sin_table(402) <= 592;
  sin_table(403) <= 593;
  sin_table(404) <= 594;
  sin_table(405) <= 595;
  sin_table(406) <= 597;
  sin_table(407) <= 598;
  sin_table(408) <= 599;
  sin_table(409) <= 601;
  sin_table(410) <= 602;
  sin_table(411) <= 603;
  sin_table(412) <= 604;
  sin_table(413) <= 606;
  sin_table(414) <= 607;
  sin_table(415) <= 608;
  sin_table(416) <= 609;
  sin_table(417) <= 611;
  sin_table(418) <= 612;
  sin_table(419) <= 613;
  sin_table(420) <= 614;
  sin_table(421) <= 616;
  sin_table(422) <= 617;
  sin_table(423) <= 618;
  sin_table(424) <= 619;
  sin_table(425) <= 621;
  sin_table(426) <= 622;
  sin_table(427) <= 623;
  sin_table(428) <= 624;
  sin_table(429) <= 626;
  sin_table(430) <= 627;
  sin_table(431) <= 628;
  sin_table(432) <= 629;
  sin_table(433) <= 631;
  sin_table(434) <= 632;
  sin_table(435) <= 633;
  sin_table(436) <= 634;
  sin_table(437) <= 636;
  sin_table(438) <= 637;
  sin_table(439) <= 638;
  sin_table(440) <= 639;
  sin_table(441) <= 640;
  sin_table(442) <= 642;
  sin_table(443) <= 643;
  sin_table(444) <= 644;
  sin_table(445) <= 645;
  sin_table(446) <= 647;
  sin_table(447) <= 648;
  sin_table(448) <= 649;
  sin_table(449) <= 650;
  sin_table(450) <= 651;
  sin_table(451) <= 653;
  sin_table(452) <= 654;
  sin_table(453) <= 655;
  sin_table(454) <= 656;
  sin_table(455) <= 657;
  sin_table(456) <= 659;
  sin_table(457) <= 660;
  sin_table(458) <= 661;
  sin_table(459) <= 662;
  sin_table(460) <= 663;
  sin_table(461) <= 665;
  sin_table(462) <= 666;
  sin_table(463) <= 667;
  sin_table(464) <= 668;
  sin_table(465) <= 669;
  sin_table(466) <= 671;
  sin_table(467) <= 672;
  sin_table(468) <= 673;
  sin_table(469) <= 674;
  sin_table(470) <= 675;
  sin_table(471) <= 676;
  sin_table(472) <= 678;
  sin_table(473) <= 679;
  sin_table(474) <= 680;
  sin_table(475) <= 681;
  sin_table(476) <= 682;
  sin_table(477) <= 684;
  sin_table(478) <= 685;
  sin_table(479) <= 686;
  sin_table(480) <= 687;
  sin_table(481) <= 688;
  sin_table(482) <= 689;
  sin_table(483) <= 690;
  sin_table(484) <= 692;
  sin_table(485) <= 693;
  sin_table(486) <= 694;
  sin_table(487) <= 695;
  sin_table(488) <= 696;
  sin_table(489) <= 697;
  sin_table(490) <= 699;
  sin_table(491) <= 700;
  sin_table(492) <= 701;
  sin_table(493) <= 702;
  sin_table(494) <= 703;
  sin_table(495) <= 704;
  sin_table(496) <= 705;
  sin_table(497) <= 707;
  sin_table(498) <= 708;
  sin_table(499) <= 709;
  sin_table(500) <= 710;
  sin_table(501) <= 711;
  sin_table(502) <= 712;
  sin_table(503) <= 713;
  sin_table(504) <= 714;
  sin_table(505) <= 716;
  sin_table(506) <= 717;
  sin_table(507) <= 718;
  sin_table(508) <= 719;
  sin_table(509) <= 720;
  sin_table(510) <= 721;
  sin_table(511) <= 722;
  sin_table(512) <= 723;
  sin_table(513) <= 724;
  sin_table(514) <= 726;
  sin_table(515) <= 727;
  sin_table(516) <= 728;
  sin_table(517) <= 729;
  sin_table(518) <= 730;
  sin_table(519) <= 731;
  sin_table(520) <= 732;
  sin_table(521) <= 733;
  sin_table(522) <= 734;
  sin_table(523) <= 735;
  sin_table(524) <= 737;
  sin_table(525) <= 738;
  sin_table(526) <= 739;
  sin_table(527) <= 740;
  sin_table(528) <= 741;
  sin_table(529) <= 742;
  sin_table(530) <= 743;
  sin_table(531) <= 744;
  sin_table(532) <= 745;
  sin_table(533) <= 746;
  sin_table(534) <= 747;
  sin_table(535) <= 748;
  sin_table(536) <= 750;
  sin_table(537) <= 751;
  sin_table(538) <= 752;
  sin_table(539) <= 753;
  sin_table(540) <= 754;
  sin_table(541) <= 755;
  sin_table(542) <= 756;
  sin_table(543) <= 757;
  sin_table(544) <= 758;
  sin_table(545) <= 759;
  sin_table(546) <= 760;
  sin_table(547) <= 761;
  sin_table(548) <= 762;
  sin_table(549) <= 763;
  sin_table(550) <= 764;
  sin_table(551) <= 765;
  sin_table(552) <= 766;
  sin_table(553) <= 767;
  sin_table(554) <= 768;
  sin_table(555) <= 769;
  sin_table(556) <= 771;
  sin_table(557) <= 772;
  sin_table(558) <= 773;
  sin_table(559) <= 774;
  sin_table(560) <= 775;
  sin_table(561) <= 776;
  sin_table(562) <= 777;
  sin_table(563) <= 778;
  sin_table(564) <= 779;
  sin_table(565) <= 780;
  sin_table(566) <= 781;
  sin_table(567) <= 782;
  sin_table(568) <= 783;
  sin_table(569) <= 784;
  sin_table(570) <= 785;
  sin_table(571) <= 786;
  sin_table(572) <= 787;
  sin_table(573) <= 788;
  sin_table(574) <= 789;
  sin_table(575) <= 790;
  sin_table(576) <= 791;
  sin_table(577) <= 792;
  sin_table(578) <= 793;
  sin_table(579) <= 794;
  sin_table(580) <= 795;
  sin_table(581) <= 796;
  sin_table(582) <= 797;
  sin_table(583) <= 798;
  sin_table(584) <= 799;
  sin_table(585) <= 800;
  sin_table(586) <= 801;
  sin_table(587) <= 802;
  sin_table(588) <= 803;
  sin_table(589) <= 804;
  sin_table(590) <= 805;
  sin_table(591) <= 806;
  sin_table(592) <= 806;
  sin_table(593) <= 807;
  sin_table(594) <= 808;
  sin_table(595) <= 809;
  sin_table(596) <= 810;
  sin_table(597) <= 811;
  sin_table(598) <= 812;
  sin_table(599) <= 813;
  sin_table(600) <= 814;
  sin_table(601) <= 815;
  sin_table(602) <= 816;
  sin_table(603) <= 817;
  sin_table(604) <= 818;
  sin_table(605) <= 819;
  sin_table(606) <= 820;
  sin_table(607) <= 821;
  sin_table(608) <= 822;
  sin_table(609) <= 823;
  sin_table(610) <= 824;
  sin_table(611) <= 824;
  sin_table(612) <= 825;
  sin_table(613) <= 826;
  sin_table(614) <= 827;
  sin_table(615) <= 828;
  sin_table(616) <= 829;
  sin_table(617) <= 830;
  sin_table(618) <= 831;
  sin_table(619) <= 832;
  sin_table(620) <= 833;
  sin_table(621) <= 834;
  sin_table(622) <= 835;
  sin_table(623) <= 835;
  sin_table(624) <= 836;
  sin_table(625) <= 837;
  sin_table(626) <= 838;
  sin_table(627) <= 839;
  sin_table(628) <= 840;
  sin_table(629) <= 841;
  sin_table(630) <= 842;
  sin_table(631) <= 843;
  sin_table(632) <= 844;
  sin_table(633) <= 844;
  sin_table(634) <= 845;
  sin_table(635) <= 846;
  sin_table(636) <= 847;
  sin_table(637) <= 848;
  sin_table(638) <= 849;
  sin_table(639) <= 850;
  sin_table(640) <= 851;
  sin_table(641) <= 851;
  sin_table(642) <= 852;
  sin_table(643) <= 853;
  sin_table(644) <= 854;
  sin_table(645) <= 855;
  sin_table(646) <= 856;
  sin_table(647) <= 857;
  sin_table(648) <= 858;
  sin_table(649) <= 858;
  sin_table(650) <= 859;
  sin_table(651) <= 860;
  sin_table(652) <= 861;
  sin_table(653) <= 862;
  sin_table(654) <= 863;
  sin_table(655) <= 863;
  sin_table(656) <= 864;
  sin_table(657) <= 865;
  sin_table(658) <= 866;
  sin_table(659) <= 867;
  sin_table(660) <= 868;
  sin_table(661) <= 868;
  sin_table(662) <= 869;
  sin_table(663) <= 870;
  sin_table(664) <= 871;
  sin_table(665) <= 872;
  sin_table(666) <= 873;
  sin_table(667) <= 873;
  sin_table(668) <= 874;
  sin_table(669) <= 875;
  sin_table(670) <= 876;
  sin_table(671) <= 877;
  sin_table(672) <= 877;
  sin_table(673) <= 878;
  sin_table(674) <= 879;
  sin_table(675) <= 880;
  sin_table(676) <= 881;
  sin_table(677) <= 881;
  sin_table(678) <= 882;
  sin_table(679) <= 883;
  sin_table(680) <= 884;
  sin_table(681) <= 885;
  sin_table(682) <= 885;
  sin_table(683) <= 886;
  sin_table(684) <= 887;
  sin_table(685) <= 888;
  sin_table(686) <= 889;
  sin_table(687) <= 889;
  sin_table(688) <= 890;
  sin_table(689) <= 891;
  sin_table(690) <= 892;
  sin_table(691) <= 892;
  sin_table(692) <= 893;
  sin_table(693) <= 894;
  sin_table(694) <= 895;
  sin_table(695) <= 895;
  sin_table(696) <= 896;
  sin_table(697) <= 897;
  sin_table(698) <= 898;
  sin_table(699) <= 898;
  sin_table(700) <= 899;
  sin_table(701) <= 900;
  sin_table(702) <= 901;
  sin_table(703) <= 901;
  sin_table(704) <= 902;
  sin_table(705) <= 903;
  sin_table(706) <= 904;
  sin_table(707) <= 904;
  sin_table(708) <= 905;
  sin_table(709) <= 906;
  sin_table(710) <= 907;
  sin_table(711) <= 907;
  sin_table(712) <= 908;
  sin_table(713) <= 909;
  sin_table(714) <= 909;
  sin_table(715) <= 910;
  sin_table(716) <= 911;
  sin_table(717) <= 912;
  sin_table(718) <= 912;
  sin_table(719) <= 913;
  sin_table(720) <= 914;
  sin_table(721) <= 914;
  sin_table(722) <= 915;
  sin_table(723) <= 916;
  sin_table(724) <= 917;
  sin_table(725) <= 917;
  sin_table(726) <= 918;
  sin_table(727) <= 919;
  sin_table(728) <= 919;
  sin_table(729) <= 920;
  sin_table(730) <= 921;
  sin_table(731) <= 921;
  sin_table(732) <= 922;
  sin_table(733) <= 923;
  sin_table(734) <= 923;
  sin_table(735) <= 924;
  sin_table(736) <= 925;
  sin_table(737) <= 925;
  sin_table(738) <= 926;
  sin_table(739) <= 927;
  sin_table(740) <= 927;
  sin_table(741) <= 928;
  sin_table(742) <= 929;
  sin_table(743) <= 929;
  sin_table(744) <= 930;
  sin_table(745) <= 931;
  sin_table(746) <= 931;
  sin_table(747) <= 932;
  sin_table(748) <= 933;
  sin_table(749) <= 933;
  sin_table(750) <= 934;
  sin_table(751) <= 935;
  sin_table(752) <= 935;
  sin_table(753) <= 936;
  sin_table(754) <= 937;
  sin_table(755) <= 937;
  sin_table(756) <= 938;
  sin_table(757) <= 938;
  sin_table(758) <= 939;
  sin_table(759) <= 940;
  sin_table(760) <= 940;
  sin_table(761) <= 941;
  sin_table(762) <= 941;
  sin_table(763) <= 942;
  sin_table(764) <= 943;
  sin_table(765) <= 943;
  sin_table(766) <= 944;
  sin_table(767) <= 945;
  sin_table(768) <= 945;
  sin_table(769) <= 946;
  sin_table(770) <= 946;
  sin_table(771) <= 947;
  sin_table(772) <= 948;
  sin_table(773) <= 948;
  sin_table(774) <= 949;
  sin_table(775) <= 949;
  sin_table(776) <= 950;
  sin_table(777) <= 950;
  sin_table(778) <= 951;
  sin_table(779) <= 952;
  sin_table(780) <= 952;
  sin_table(781) <= 953;
  sin_table(782) <= 953;
  sin_table(783) <= 954;
  sin_table(784) <= 954;
  sin_table(785) <= 955;
  sin_table(786) <= 956;
  sin_table(787) <= 956;
  sin_table(788) <= 957;
  sin_table(789) <= 957;
  sin_table(790) <= 958;
  sin_table(791) <= 958;
  sin_table(792) <= 959;
  sin_table(793) <= 959;
  sin_table(794) <= 960;
  sin_table(795) <= 961;
  sin_table(796) <= 961;
  sin_table(797) <= 962;
  sin_table(798) <= 962;
  sin_table(799) <= 963;
  sin_table(800) <= 963;
  sin_table(801) <= 964;
  sin_table(802) <= 964;
  sin_table(803) <= 965;
  sin_table(804) <= 965;
  sin_table(805) <= 966;
  sin_table(806) <= 966;
  sin_table(807) <= 967;
  sin_table(808) <= 967;
  sin_table(809) <= 968;
  sin_table(810) <= 968;
  sin_table(811) <= 969;
  sin_table(812) <= 969;
  sin_table(813) <= 970;
  sin_table(814) <= 970;
  sin_table(815) <= 971;
  sin_table(816) <= 971;
  sin_table(817) <= 972;
  sin_table(818) <= 972;
  sin_table(819) <= 973;
  sin_table(820) <= 973;
  sin_table(821) <= 974;
  sin_table(822) <= 974;
  sin_table(823) <= 975;
  sin_table(824) <= 975;
  sin_table(825) <= 976;
  sin_table(826) <= 976;
  sin_table(827) <= 977;
  sin_table(828) <= 977;
  sin_table(829) <= 978;
  sin_table(830) <= 978;
  sin_table(831) <= 978;
  sin_table(832) <= 979;
  sin_table(833) <= 979;
  sin_table(834) <= 980;
  sin_table(835) <= 980;
  sin_table(836) <= 981;
  sin_table(837) <= 981;
  sin_table(838) <= 982;
  sin_table(839) <= 982;
  sin_table(840) <= 983;
  sin_table(841) <= 983;
  sin_table(842) <= 983;
  sin_table(843) <= 984;
  sin_table(844) <= 984;
  sin_table(845) <= 985;
  sin_table(846) <= 985;
  sin_table(847) <= 986;
  sin_table(848) <= 986;
  sin_table(849) <= 986;
  sin_table(850) <= 987;
  sin_table(851) <= 987;
  sin_table(852) <= 988;
  sin_table(853) <= 988;
  sin_table(854) <= 988;
  sin_table(855) <= 989;
  sin_table(856) <= 989;
  sin_table(857) <= 990;
  sin_table(858) <= 990;
  sin_table(859) <= 990;
  sin_table(860) <= 991;
  sin_table(861) <= 991;
  sin_table(862) <= 992;
  sin_table(863) <= 992;
  sin_table(864) <= 992;
  sin_table(865) <= 993;
  sin_table(866) <= 993;
  sin_table(867) <= 993;
  sin_table(868) <= 994;
  sin_table(869) <= 994;
  sin_table(870) <= 995;
  sin_table(871) <= 995;
  sin_table(872) <= 995;
  sin_table(873) <= 996;
  sin_table(874) <= 996;
  sin_table(875) <= 996;
  sin_table(876) <= 997;
  sin_table(877) <= 997;
  sin_table(878) <= 997;
  sin_table(879) <= 998;
  sin_table(880) <= 998;
  sin_table(881) <= 998;
  sin_table(882) <= 999;
  sin_table(883) <= 999;
  sin_table(884) <= 999;
  sin_table(885) <= 1000;
  sin_table(886) <= 1000;
  sin_table(887) <= 1000;
  sin_table(888) <= 1001;
  sin_table(889) <= 1001;
  sin_table(890) <= 1001;
  sin_table(891) <= 1002;
  sin_table(892) <= 1002;
  sin_table(893) <= 1002;
  sin_table(894) <= 1003;
  sin_table(895) <= 1003;
  sin_table(896) <= 1003;
  sin_table(897) <= 1004;
  sin_table(898) <= 1004;
  sin_table(899) <= 1004;
  sin_table(900) <= 1005;
  sin_table(901) <= 1005;
  sin_table(902) <= 1005;
  sin_table(903) <= 1005;
  sin_table(904) <= 1006;
  sin_table(905) <= 1006;
  sin_table(906) <= 1006;
  sin_table(907) <= 1007;
  sin_table(908) <= 1007;
  sin_table(909) <= 1007;
  sin_table(910) <= 1007;
  sin_table(911) <= 1008;
  sin_table(912) <= 1008;
  sin_table(913) <= 1008;
  sin_table(914) <= 1008;
  sin_table(915) <= 1009;
  sin_table(916) <= 1009;
  sin_table(917) <= 1009;
  sin_table(918) <= 1010;
  sin_table(919) <= 1010;
  sin_table(920) <= 1010;
  sin_table(921) <= 1010;
  sin_table(922) <= 1011;
  sin_table(923) <= 1011;
  sin_table(924) <= 1011;
  sin_table(925) <= 1011;
  sin_table(926) <= 1011;
  sin_table(927) <= 1012;
  sin_table(928) <= 1012;
  sin_table(929) <= 1012;
  sin_table(930) <= 1012;
  sin_table(931) <= 1013;
  sin_table(932) <= 1013;
  sin_table(933) <= 1013;
  sin_table(934) <= 1013;
  sin_table(935) <= 1013;
  sin_table(936) <= 1014;
  sin_table(937) <= 1014;
  sin_table(938) <= 1014;
  sin_table(939) <= 1014;
  sin_table(940) <= 1015;
  sin_table(941) <= 1015;
  sin_table(942) <= 1015;
  sin_table(943) <= 1015;
  sin_table(944) <= 1015;
  sin_table(945) <= 1015;
  sin_table(946) <= 1016;
  sin_table(947) <= 1016;
  sin_table(948) <= 1016;
  sin_table(949) <= 1016;
  sin_table(950) <= 1016;
  sin_table(951) <= 1017;
  sin_table(952) <= 1017;
  sin_table(953) <= 1017;
  sin_table(954) <= 1017;
  sin_table(955) <= 1017;
  sin_table(956) <= 1017;
  sin_table(957) <= 1018;
  sin_table(958) <= 1018;
  sin_table(959) <= 1018;
  sin_table(960) <= 1018;
  sin_table(961) <= 1018;
  sin_table(962) <= 1018;
  sin_table(963) <= 1019;
  sin_table(964) <= 1019;
  sin_table(965) <= 1019;
  sin_table(966) <= 1019;
  sin_table(967) <= 1019;
  sin_table(968) <= 1019;
  sin_table(969) <= 1019;
  sin_table(970) <= 1019;
  sin_table(971) <= 1020;
  sin_table(972) <= 1020;
  sin_table(973) <= 1020;
  sin_table(974) <= 1020;
  sin_table(975) <= 1020;
  sin_table(976) <= 1020;
  sin_table(977) <= 1020;
  sin_table(978) <= 1020;
  sin_table(979) <= 1021;
  sin_table(980) <= 1021;
  sin_table(981) <= 1021;
  sin_table(982) <= 1021;
  sin_table(983) <= 1021;
  sin_table(984) <= 1021;
  sin_table(985) <= 1021;
  sin_table(986) <= 1021;
  sin_table(987) <= 1021;
  sin_table(988) <= 1021;
  sin_table(989) <= 1022;
  sin_table(990) <= 1022;
  sin_table(991) <= 1022;
  sin_table(992) <= 1022;
  sin_table(993) <= 1022;
  sin_table(994) <= 1022;
  sin_table(995) <= 1022;
  sin_table(996) <= 1022;
  sin_table(997) <= 1022;
  sin_table(998) <= 1022;
  sin_table(999) <= 1022;
  sin_table(1000) <= 1022;
  sin_table(1001) <= 1022;
  sin_table(1002) <= 1022;
  sin_table(1003) <= 1022;
  sin_table(1004) <= 1023;
  sin_table(1005) <= 1023;
  sin_table(1006) <= 1023;
  sin_table(1007) <= 1023;
  sin_table(1008) <= 1023;
  sin_table(1009) <= 1023;
  sin_table(1010) <= 1023;
  sin_table(1011) <= 1023;
  sin_table(1012) <= 1023;
  sin_table(1013) <= 1023;
  sin_table(1014) <= 1023;
  sin_table(1015) <= 1023;
  sin_table(1016) <= 1023;
  sin_table(1017) <= 1023;
  sin_table(1018) <= 1023;
  sin_table(1019) <= 1023;
  sin_table(1020) <= 1023;
  sin_table(1021) <= 1023;
  sin_table(1022) <= 1023;
  sin_table(1023) <= 1023;

  addr_tmp <= conv_integer(unsigned(addr_i));
  sin_tmp  <= conv_std_logic_vector(sin_table(addr_tmp),10);
  
  sin_o    <= sin_tmp;

end rtl;
