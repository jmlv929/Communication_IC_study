
--============================================================================--
--                                   ARCHITECTURE                             --
--============================================================================--

architecture RTL of aes_subbytes is

--------------------------------------------------------------- Type declaration
type s_box_type   is array (255 downto 0) of std_logic_vector (7 downto 0);
-------------------------------------------------------- End of Type declaration

-------------------------------------------------------------- S-Box declaration
-- These are the values in the S-Box used to make the State transformation:
constant s_box_ct : s_box_type
          := ("00010110", "10111011", "01010100", "10110000", -- 16, BB, 54, B0.
              "00001111", "00101101", "10011001", "01000001", -- 0F, 2D, 99, 41.
              "01101000", "01000010", "11100110", "10111111", -- 68, 42, E6, BF.
              "00001101", "10001001", "10100001", "10001100", -- 0D, 89, A1, 8C.

              "11011111", "00101000", "01010101", "11001110", -- DF, 28, 55, CE.
              "11101001", "10000111", "00011110", "10011011", -- E9, 87, 1E, 9B.
              "10010100", "10001110", "11011001", "01101001", -- 94, 8E, D9, 69.
              "00010001", "10011000", "11111000", "11100001", -- 11, 98, F8, E1.

              "10011110", "00011101", "11000001", "10000110", -- 9E, 1D, C1, 86.
              "10111001", "01010111", "00110101", "01100001", -- B9, 57, 35, 61.
              "00001110", "11110110", "00000011", "01001000", -- 0E, F6, 03, 48.
              "01100110", "10110101", "00111110", "01110000", -- 66, B5, 3E, 70.

              "10001010", "10001011", "10111101", "01001011", -- 8A, 8B, BD, 4B.
              "00011111", "01110100", "11011101", "11101000", -- 1F, 74, DD, E8.
              "11000110", "10110100", "10100110", "00011100", -- C6, B4, A6, 1C.
              "00101110", "00100101", "01111000", "10111010", -- 2E, 25, 78, BA.

              "00001000", "10101110", "01111010", "01100101", -- 08, AE, 7A, 65.
              "11101010", "11110100", "01010110", "01101100", -- EA, F4, 56, 6C.
              "10101001", "01001110", "11010101", "10001101", -- A9, 4E, D5, 8D.
              "01101101", "00110111", "11001000", "11100111", -- 6D, 37, C8, E7.

              "01111001", "11100100", "10010101", "10010001", -- 79, E4, 95, 91.
              "01100010", "10101100", "11010011", "11000010", -- 62, AC, D3, C2.
              "01011100", "00100100", "00000110", "01001001", -- 5C, 24, 06, 49.
              "00001010", "00111010", "00110010", "11100000", -- 0A, 3A, 32, E0.

              "11011011", "00001011", "01011110", "11011110", -- DB, 0B, 5E, DE,
              "00010100", "10111000", "11101110", "01000110", -- 14, B8, EE, 46.
              "10001000", "10010000", "00101010", "00100010", -- 88, 90, 2A, 22.
              "11011100", "01001111", "10000001", "01100000", -- DC, 4F, 81, 60.

              "01110011", "00011001", "01011101", "01100100", -- 73, 19, 5D, 64.
              "00111101", "01111110", "10100111", "11000100", -- 3D, 7E, A7, C4.
              "00010111", "01000100", "10010111", "01011111", -- 17, 44, 97, 5F.
              "11101100", "00010011", "00001100", "11001101", -- EC, 13, 0C, CD.

              "11010010", "11110011", "11111111", "00010000", -- D2, F3, FF, 10.
              "00100001", "11011010", "10110110", "10111100", -- 21, DA, B6, BC.
              "11110101", "00111000", "10011101", "10010010", -- F5, 38, 9D, 92.
              "10001111", "01000000", "10100011", "01010001", -- 8F, 40, A3, 51.

              "10101000", "10011111", "00111100", "01010000", -- A8, 9F, 3C, 50.
              "01111111", "00000010", "11111001", "01000101", -- 7F, 02, F9, 45.
              "10000101", "00110011", "01001101", "01000011", -- 85, 33, 4D, 43.
              "11111011", "10101010", "11101111", "11010000", -- FB, AA, EF, D0.

              "11001111", "01011000", "01001100", "01001010", -- CF, 58, 4C, 4A.
              "00111001", "10111110", "11001011", "01101010", -- 39, BE, CB, 6A.
              "01011011", "10110001", "11111100", "00100000", -- 5B, B1, FC, 20.
              "11101101", "00000000", "11010001", "01010011", -- ED, 00, D1, 53.

              "10000100", "00101111", "11100011", "00101001", -- 84, 2F, E3, 29.
              "10110011", "11010110", "00111011", "01010010", -- B3, D6, 3B, 52.
              "10100000", "01011010", "01101110", "00011011", -- A0, 5A, 6E, 1B.
              "00011010", "00101100", "10000011", "00001001", -- 1A, 2C, 83, 09.

              "01110101", "10110010", "00100111", "11101011", -- 75, B2, 27, EB.
              "11100010", "10000000", "00010010", "00000111", -- E2, 80, 12, 07.
              "10011010", "00000101", "10010110", "00011000", -- 9A, 05, 96, 18.
              "11000011", "00100011", "11000111", "00000100", -- C3, 23, C7, 04.

              "00010101", "00110001", "11011000", "01110001", -- 15, 31, D8, 71.
              "11110001", "11100101", "10100101", "00110100", -- F1, E5, A5, 34.
              "11001100", "11110111", "00111111", "00110110", -- CC, F7, 3F, 36.
              "00100110", "10010011", "11111101", "10110111", -- 26, 93, FD, B7.

              "11000000", "01110010", "10100100", "10011100", -- C0, 72, A4, 9C.
              "10101111", "10100010", "11010100", "10101101", -- AF, A2, D4, AD.
              "11110000", "01000111", "01011001", "11111010", -- F0, 47, 59, FA.
              "01111101", "11001001", "10000010", "11001010", -- 7D, C9, 82, CA.

              "01110110", "10101011", "11010111", "11111110", -- 76, AB, D7, FE.
              "00101011", "01100111", "00000001", "00110000", -- 2B, 67, 01, 30.
              "11000101", "01101111", "01101011", "11110010", -- C5, 6F, 6B, F2.
              "01111011", "01110111", "01111100", "01100011");-- 7B, 77, 7C, 63.
------------------------------------------------------- End of S-Box declaration

------------------------------------------------------------- Signal declaration
signal byte_in0  : std_logic_vector (7 downto 0);
signal byte_in1  : std_logic_vector (7 downto 0);
signal byte_in2  : std_logic_vector (7 downto 0);
signal byte_in3  : std_logic_vector (7 downto 0);
signal byte_out0 : std_logic_vector (7 downto 0);
signal byte_out1 : std_logic_vector (7 downto 0);
signal byte_out2 : std_logic_vector (7 downto 0);
signal byte_out3 : std_logic_vector (7 downto 0);
------------------------------------------------------ End of signal declaration

begin

  ---------------------------------------------------------- Byte transformation
  -- This block transforms the 32-bit input lines into 8-bits signals and the
  -- result into 32-bit output lines.
  byte_in0 <= word_in ( 7 downto  0);
  byte_in1 <= word_in (15 downto  8);
  byte_in2 <= word_in (23 downto 16);
  byte_in3 <= word_in (31 downto 24);
  word_out <= byte_out3 & byte_out2 & byte_out1 & byte_out0;
  --------------------------------------------------- End of Byte transformation

  -------------------------------------------------------- Column Transformation
  -- This process calculates the transformations that correspond to each byte
  -- in one of the matrix column. The calculation is done looking at the
  -- corresponding value in the S-Box.
  byte_out0 <= s_box_ct (conv_integer (byte_in0));
  byte_out1 <= s_box_ct (conv_integer (byte_in1));
  byte_out2 <= s_box_ct (conv_integer (byte_in2));
  byte_out3 <= s_box_ct (conv_integer (byte_in3));
  ------------------------------------------------- End of Column Transformation

end RTL;
