
--------------------------------------------------------------------------------
-- Architecture
--------------------------------------------------------------------------------
architecture rtl of ha is

begin  -- rtl

  c <= x and y;
  s <= x xor y;

end rtl;
