
--------------------------------------------------------------------------------
-- End of file
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--       ------------      Project : WiLD
--    ,' GoodLuck ,'      RCSfile: sine_table_rom_pkg.vhd,v   
--   '-----------'     Author: DR \*
--
--  Revision: 1.1   
--  Date: 1999.12.31
--  State: Exp  
--  Locker:   
--------------------------------------------------------------------------------
--
-- Description : Package for sine_table_rom.
--
--------------------------------------------------------------------------------
--
--  Source: ./git/COMMON/IPs/WILD/MODEM802_11a2/sine_table_rom/vhdl/rtl/sine_table_rom_pkg.vhd,v  
--  Log: sine_table_rom_pkg.vhd,v  
-- Revision 1.1  2003/03/13 15:26:20  Dr.A
-- Initial revision
--
--
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
-- Library
--------------------------------------------------------------------------------
library IEEE; 
    use IEEE.STD_LOGIC_1164.ALL; 

--------------------------------------------------------------------------------
-- Package
--------------------------------------------------------------------------------
package sine_table_rom_pkg is


--------------------------------------------------------------------------------
-- Components list declaration done by <fb> script.
--------------------------------------------------------------------------------
----------------------
-- File: sine_table_rom.vhd
----------------------
  component sine_table_rom
  port (
     addr_i   : in  std_logic_vector(9 downto 0); -- input angle
     sin_o    : out std_logic_vector(9 downto 0)  -- output sine
  );

  end component;



 
end sine_table_rom_pkg;
