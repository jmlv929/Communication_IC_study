

--------------------------------------------------------------------------------
-- Architecture
--------------------------------------------------------------------------------
architecture RTL of kalman_lut is

  ------------------------------------------------------------------------------
  -- Types
  ------------------------------------------------------------------------------

  ------------------------------------------------------------------------------
  -- Signals
  ------------------------------------------------------------------------------
  signal k_int  : natural range 1 to 247;
  signal km_int : natural range 777 to 1023;

--------------------------------------------------------------------------------
-- Architecture Body
--------------------------------------------------------------------------------
begin

  with k_index select
    k_int <=
    247 when "000000",
    199 when "000001",
      1 when "000010",
    171 when "000011",
    156 when "000100",
    142 when "000101",
    129 when "000110",
    118 when "000111",
    107 when "001000",
     98 when "001001",
     89 when "001010",
     81 when "001011",
     74 when "001100",
     67 when "001101",
     61 when "001110",
     56 when "001111",
     51 when "010000",
     46 when "010001",
     42 when "010010",
     39 when "010011",
     35 when "010100",
     32 when "010101",
     29 when "010110",
     27 when "010111",
     24 when "011000",
     22 when "011001",
     20 when "011010",
     18 when "011011",
     17 when "011100",
     15 when "011101",
     14 when "011110",
     13 when "011111",
     12 when "100000",
     10 when "100001",
     10 when "100010",
      9 when "100011",
      8 when "100100",
      7 when "100101",
      7 when "100110",
      6 when "100111",
      5 when "101000",
      5 when "101001",
      5 when "101010",
      4 when "101011",
      4 when "101100",
      3 when "101101",
      3 when "101110",
      3 when "101111",
      3 when "110000",
      2 when "110001",
      2 when "110010",
      2 when "110011",
      2 when "110100",
      2 when "110101",
      1 when "110110",
      1 when "110111",
      1 when "111000",
      1 when "111001",
      1 when "111010",
      1 when "111011",
      1 when "111100",
      1 when "111101",
      1 when "111110",
      1 when "111111",
      1 when others;   



  with k_index select
    km_int <=
     777 when "000000",
     825 when "000001",
    1023 when "000010",
     853 when "000011",
     868 when "000100",
     882 when "000101",
     895 when "000110",
     906 when "000111",
     917 when "001000",
     926 when "001001",
     935 when "001010",
     943 when "001011",
     950 when "001100",
     957 when "001101",
     963 when "001110",
     968 when "001111",
     973 when "010000",
     978 when "010001",
     982 when "010010",
     985 when "010011",
     989 when "010100",
     992 when "010101",
     995 when "010110",
     997 when "010111",
    1000 when "011000",
    1002 when "011001",
    1004 when "011010",
    1006 when "011011",
    1007 when "011100",
    1009 when "011101",
    1010 when "011110",
    1011 when "011111",
    1012 when "100000",
    1014 when "100001",
    1014 when "100010",
    1015 when "100011",
    1016 when "100100",
    1017 when "100101",
    1017 when "100110",
    1018 when "100111",
    1019 when "101000",
    1019 when "101001",
    1019 when "101010",
    1020 when "101011",
    1020 when "101100",
    1021 when "101101",
    1021 when "101110",
    1021 when "101111",
    1021 when "110000",
    1022 when "110001",
    1022 when "110010",
    1022 when "110011",
    1022 when "110100",
    1022 when "110101",
    1023 when "110110",
    1023 when "110111",
    1023 when "111000",
    1023 when "111001",
    1023 when "111010",
    1023 when "111011",
    1023 when "111100",
    1023 when "111101",
    1023 when "111110",
    1023 when "111111",
    1023 when others;

  k_o  <= conv_std_logic_vector(k_int, 10);
  km_o <= conv_std_logic_vector(km_int, 10);
  
end RTL;
